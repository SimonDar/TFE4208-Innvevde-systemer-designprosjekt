��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j0y�ߞ��'DmP"l�8Ws����3#�P����P�ɻ��v�B�*����ހٗ��l�I�$JE�����X�(�>���'v���)U:���si����mY��������f}���/ p�2P�W���v�R�9d��$h�E�o���kI���c�z%�y��	E<|���Ur��~����M��`(���)dDP�>��B� G���^E�<.���t`
��0�ڙv���I�KH߀ܚV��!�
�!֑|�f���#G&Q��%���َ!}�?ғ�H�
�?�{1�,�w�JG}CtVa���+�tl �P_G:���E�v�E$b�S�����0�@!�ʁ::�� �y'��wp��Ú��Jk`�14���VbIO����֪J��[�Bi�k·�h
���j_R�-����&�׍�m��9�Ϸy(\7A'ޏ�}	҈(���)��2j8���5)vLP���b��z?��Ѣ"�/���b�@�V������fY�:]>��bN�<=�3m�7��M\NP"���j1S�{ن�r�A���et�«���Y��sW?K	L���C�ypnk\.��L/�l�ћ�X5�oѪO���/&�;%��2��`�ě��j}6�8/m^@�D��KB�%/
�������pRa��PF�4�
ݔ#Z�*W0�@;2+�{�$ri�`]���HCE���l�����P�;}��uM����B��f�k%V���Ly'���
O���ʮ�h�0����|4OԢ+�}�$�t��faC�C��ܞ��ޒ�����A������҅ӱ	H�ul�Ɉ\�<R��V��WgA�I!/����^x�Ra0[F�N7om�K_E�A���z?e�ր�@�G�
�A�8�i�"���'��9{i���R�HR�y��Yp�䝔6�c$��@�d��;#�n��.�A��{ިǫ�I�L<��[8�,w�)�����'�: �ߑ�1�	c-���*������U���~�o�6���UO���#ޝ>��#GiG&&���Ήy�*���AR�|L�Bl/�5��R�]Kh�f�i6n��G�}ds�vbW�ha�)d��ݪ~�*n�|4zֈ��������r��>��Qh?EY�?��w
_��T�j�坸��������8ܖy��8ۅ�ѣ�+��­���2/B��
�E�jK�O��ǧ� (ȟ��h0JGm��;��`�~����],6��	����o�ԑ�T&�����UG�w����?M�C�q�Bw�2�!O_����_-тG�;�c�r�-y�'�Yi����*ޘ���U)b�_���@�~CKuz�,�hF^���S�х2XUv�I��!&/��h!%G5��.��R�r�d,�mP)g~���{Qt����tC�s�0��5 ���F�ar�ˮ���H��o�ם����`T2&fO)�~�p��2��ʨ�`SYi#"���J��/	��r��9[#ζ��y�^��ԅ
�)�6AO��Dz��*o�����ŒB�1�by��R����(����}��� =B�P���M�o-�nf[)^X4�,����)u$��8��BSٵXcHZE�~���ܾW�iL��OLK`����Q�Q�ݸ���k��R7���y`J��M�Ǎ�#4K7{\ ��р��Aw��/�����0�SU(1��@�DA0�����C��)��Q��9;�:���΅-#� a����@%�a�j���y�vhNRX�=��^�w?2�ŭ3���B�������a.�w��3��k�N�X��?;��$QvB�ᦊU\M%_���Sܶ5������=79E����������W
Q[��8�6ߍ�/t���}]�6Ͽ�S�{5p�y��-,��O[���Q����j�S��u���J�?��C�/��"����0�~�t��hf����6AN K�7�y�$����R�A�Όo6�#�#<]4S�	UJ�HXoR�����B�/�^d��W�|B�V��mq��|�,v�����ݞ�
&����A�k�bX��as��>W�E��7�ۆ�\�h&�Z����=Y�AA�:��R�e�����L`��Ґ��(K��o�^��P���I!^*��S�V��=�[�S�wO��8n�3�O�@e���0�c�������1@��F�vn׫�j���Ӹ-.1����
�_H������&`�뛄:��v�м��~�^���H�_��;�uS��_(Vg�lpa��*4z���K�0lS��.\+�!�4�=�lp����7|u�|���f�}�Kl��|1T��N�9?���7��0\N�zQD�7�{N�io]�L�p�ȡ���$�n 5i)��F�o�P Z�!P+�xI�K�e�C��oW��z<J�hZ��1�&b}��|�a�tg`NUY��=��~�u,~ȏ$>�j3'&$�*~9��Zk)�q���8����v���$�";_6����vg�t��N=a�ߡ�w�֙��~W'��	���������.8���d�!���a��QR��u��C�����[�%N�K�Q�p/h�In�]���P<���W:Ț�����7�^�ŭ,���������C'bX� a��A��l,�k���D�m������'��Q�@+�ɶ��EVu�S^�|�@�+0V\�Z�4�(͹������]�=l����J�}�aā�Z����}�O7F�)�� ���˲���cj�r�"G'�>�b�u'X�W������ �ޡ��"g'55���r	y��zI���m���ľO�䑕>Ĩ&��A�Ã���򱝪�N�Ҿ? y��	ʺƝ]����e�u��däB\��A6s�/u��I;�`��r�/��tfn�g.����.��8o��x�L�͡��`��e<���J����WdwA^���QÚt�>U��uS�%�B3��b��ݞ�*ǣ�L���âQ����{��{�%/(�딩H��M���2��9/=����Gy	��?�K[ ���-x?�^.��h�
�ĳ�x�e{MXO��>�A����i)zߧH-��a�r�SO���7��Z<� �ڼ����<ŝ�U�@�m��F�~�J� �Xp�� )F`9,��ְ�9�&��4wwk��/�.��k��k��2u�?8<�r���D|�l>���۷N(#��2���!�S�&�{�+��A�#�����,lob�8��(N�C��v���-|#ɠ�F��!(��� �VA��|w�����.m)��|�۳ްqn5�y�C��4YF��p2�_�\�ɴ`H} 7�u�C,_����K��8?�*#"��AR)�`�_T�c��UĿ�'x�/��N4�(�m�%�
�D	;�]2+)k0�+�dm���]�+���eo9�a�BMG=���d﷾�`Z�KD������,R��c��NɿBz++F�Uq=K:�,�X-�/[ao	�9y������m��5C��.|���]��7�td��n�}3�e[�����U���R&A!j�uA{�DM��2 �u_Ixq=���@R��'�DD�퓏wtZd_n5��_r�n�c��s��N�r!�{t�����8�u��J<���W`��Q��ϫn��h���T4ߕ�i���_C�S���9�������)�<��kU��P/����(�y��.��KR��Qka�vú8eD��fi?���֓�~�s?���٪Y�=��y��'��]յ*��	��[���(�8��Go؍E,B4w7q]�:��8��1��Ռ7�A�fF�V	�n0�5�rӢ+��3���#T58��aFѶ�O\�l̶�2��%e����WCy�2���q=�[!����
�V�j��͑J�Q^s���H�V��TDܬ�Bݳ�Z�`�T������l�q�9��R��BK