��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j0y�ߞ��'DmP"l�8Ws����3#�P����P�ɻ��v�B�*����ހٗ��l�I�$JE�����X�(�>���'v���)U:���si����mY��������f}���/ p�2P�W���v�R�9d��$h�E�o���kI���c�z%�y��	E<|���Ur��~����M��`(���)dDP�>��B� G��*�g�6u5�B����oMC����![gL� h:o��`+,jE"�+ԥL�?x�Ml;�����}�;�'K��߇F��!:�I�Y'_�J����l�%>j���qD~����1�O��T���r�v�^O�B7߮��>s5�&K��	>ɖ������:�u'i�ת��P�~Y;q=�{XS���&��[���&�~р�rI� �}Jg���Se��W����t�$bn��`r
Ė�+��=_��P�e�
k���ł;�۽Όo�p���!�|T�9�I��W7;G���~�z=A��	��_,���,�v&����8^w獽�تJ��6��-ǶDϴ�_�70!��Ҳ��_Tt�*�|:aԚ�����'c����u>�?W^�-��!���f�Sk
��e�q1u�t�B��a)]��6˰��6z|�͓2�����Px"���Bk��0�
0\����yq�*�<��6?tU� o، {u`��e��� ��=d�&��2���J��Ͱ�W����zX���,@`��N�h6V�~�E+A�~�¢M�玻E�������ī�kl���l#����1����������`�~Q����3R��'����P[�zsY3����� B>�h�, )��t��������~7�T�����NX6�j�apjs�'	���bǝ>����h���H��3�+��m��ˈW��T�{�@�?*�fq�V4���"�w9k2Z�P�q\xn�8�g�wg�Q  �a��#N��\ӏ�l�B��Lޫv�Ċku�����?��z��P��\2��%P�8���eC�6��q#�C�%�#M��9'�2O�	�%[��{@�!�H�.X��i�N��窝�8��?��R_樒����so�Q@Ap�>��=�M=7j�Љ��e�s+q��6n��AM�r\W?�G8��ǰ��jR0S_�B�!�I$�^�hj����=A3�=뙘�M@ ?��S�Ӳ���Y�_I)�yC	~��:S���r�-�)s(�D?����G��
��~;M�kc�U��q[�ld�ɫ��,��Ua�]+N���/6����S��o_�?����l 'j�v�<��hԥ����%�j|q|A�I�A`=� 3��z����f���jD�a
\��"%G>�N�B�o������M�l�lbo����ٴ��A5�m�bZu\��@���a���*	����Fe9�yǆZ�ڡ��^d��Ā������� J��2�e�������g����Rs29�q/�rC_@�k�B�g"�'�~�"PwYB���tlӪ�P����S��xʟOT��g��<:nHE�<��aI���%�f�#ӌ��ɛ5yo�zغA$��%��%�L�Z����$;7g]�!ܢk�9Hj��!���]9�����R��;�s�7?|\��<i�F
9f_��QK�J�����T�%�ph�FO4e�{���Ѹ֫�a��o�O�56
f���̖0�A��ӷ&��PD���`u\����s��&~)���n�YIF���F��ˮ	F�d���9�$[�骙�X�_���@�ρ-����n~��:�|o��*������k�P�z�wAC��iǽ��q5�):]��� ڳ+�V��9n�w�f?�ք��}���j��A��@_ d�m��-aSp�^��C0��Ě fo�.����@��R��`�:D��/�K�m�=�V���ʤ?M�.����:&��{��C���M��f`t�ﯧAc�5�(�\`t���G0Y������0vA$�DE���K��밐����'�aϢP�[@��>?A۲HPW��D<�l����cn���m�C�������N�1N�9����ue�����3n��4����Ϝ��%��͗V!ą���#�$��Ӟ�^�91g|W̗H��l�K�V�p[�(v1�%��27���?:��3��u���K�B_n�]�,H�֟)H��S��}50�bc�V|H\�����{��3/|Y�1�g���rh��nq۳·�\��|�AWq��t
I���k��e�eS��J����5A�$�A�ģ��\���4�B.�`�����|�I��l ����(�*3�5��{v2	$,��
o���cK�]A|r�{�ḅ<o��Z%�i>ܾ�[�������#�����b(���f��(�箱�.�o���*l�;�à�`����"?�r���{mIF��4��Ac�Qe����\�HDX}��q�۹T_��%q�3�b��n���,�lX.������������Q��Ck��	��	���ŀW���rBxNaP�H��e�A��q�LO��y�Lzu��Q��o���V�r��k�͐�7���Ʈ��=��`�P%���{J?�F&��{��aH���<^A�І7��f�0[��wg4�%�ke@���~HF)訡�o*�I�����Z4��Vdj'�K1=o2I�*�8#2ķ:���.�0}�(!�O�6������v]sK���Q*���Ў 1*�Uie*&:���c`�"�8k�z#H��QI�x{��۲����Y� ~~�ʛe��'��G��y9�~�mF�\R���TX{ʠ�x�J�(�������u����I�3��-Եa�-P�t8�o%	�F���y/H��;�4�,d���|��X�!�ݖ����1�$��xώϱg����}��� ����|�L��1�[-j����2�ܦ��K\�6�s�>�him�w3+(���Ǘ�CXʱT��PߧA��4�%]�C���$�����#��Q�.��u��'�t�E�G�T�Fq~�� w]�]L<�L�&"P푋i��>�s�ɢ��WD�'7�pz��:�)�Р�$����RP�����X
ɼ��M��������d�D��נV>�mrk����R�e���ƨ9�ë�ΦG_�[|��`_��b�>�M!�u�N��.�8�!ڞ�Z؀%kn{e�m{~ib'���t���Qn���m���&G��2lc��D�x���R��P���oR`[�T�x��8|���3lW�cN2�V�Ĕ �rh�V�X��-�&Ú��a�A�����~LF��<��%�로1`0�.-���p	���j��baGc_q�}�n���<9��1<"@��(���!�Vj�&69l0�z��`h������늝��QG滠u橶n��(:�'r �G�gu�5d7je�GDL�����j�G�}h�Y<g~�	~P�ǨO-G��A������lNJlB�_��q�:���ެX�{g�V��J�����s�bM~�B�W<[8b��jb�G]��R8���CD=U�-q��?�	��- ���ȓFmUQ�gSu��.����p�v1��Ŋ�d�޳If�$u�m(��L�s��Ľg�rc�n����FyI@⌮X�e���'ϨQG�x{�v&��.�bQ�M\>V�2V����y�6[�/p"U���f�I����(cS�Ld�}Pvq�'��!�C��RA��kK:���#O��0~3�EYٷ8�<�f�Ӎ�N ��S��걶�ݺv���Ўoi9�JE�� /]�zs��MB�s��Ƶ��(���PM�vx�Dn�~�5�4f��պ(3oʲ��4�c�� Wy	���Ub�����-`_�/�<�1�5,vKDp���8�Z]a
�B��
g����k��r:U�měu�Sc;�L�Y�J��đ��彥7���<^|6S/$R�-rs�3���Qjb?E4Ɓ��Pbi�u��J���3��!��Ң��� `	�u�9YAPiE]o>6�Ff<	�#�._�]��0�Ӌ��_�ZŢ����qv��/f(�V.y9="����3���M,���6.�- �=�I��~�b�kY`+�.|+޴҃�7Ps>�M��x����W�?��°{�@��]�����R��S�%�r�gqs�ش�-��鳰�V$P��׵�h��f�8�#=@H���:1e7XV�
�����&�����>����D\8K����@�����Q�j���O<>kV|�6 +�2G3�c;���@��Ld۞?���~%��l�=>�*c�{�m@B�_�7\G�#}5㵲qΖ����GR'�ݳx��8p (��?!���;&��~H� ���!t�u���6&D�j�t�h����.V��&o5�����k捷�R�7�0�E�<�< �9�vMV5O����7|�t�.%����GH��4:i�)Om05�7�ɭR�{j!@�A�O��W�𒾴;�7F�e��jֲ��'�8n�럺�e�2R��C��7_a\��l�FAWTKǡ��7 ��Z�o��"mbv*���C�H�Z�F��/`[,�����L|���So&U}�T�Ȯ�l�4�!x�,6�[��g$��z��L����d����0�x�(���"�k��{��C�e;�{�H�'M���M�x8s�=���7�7�pb-��6�\`�u�(�x�Bp}%�f���Yf������p~�au�T�[����6���&��ŕ�i���f�_K�o�;E�5��)�Wg�*��Ę���!ֺ[/)�D3_��K�r��%��k8B��z��$��B�o��N�=�<�N3�}	_��2	7������Y�W+_#�.�R	P�(���S4`${��+���ꮜA�eEh�H�ܵM{K-����x�>?s��c&8;6��ӡ�}$;׎�6�9{�:1[�l��Vz�����伀�gw|�޴ۀȷLl�1�jp��h��@I��Z֊���r�KY��7������u��mm?="�{	��W�Q}4�y��TvdF�Hdn��NImʬy���e�ᎉe���2���1��E0�u�ְ��c�����=aA��j�(��V��|�<?IhI��h�M\0�e&,,*2���7�����t�T?���<���k����+�=F=W��cD�괜�K�|4� ������(�@����%��|0�N�e��b����͊��g���w��<hT�H����3��S�_%�?Нw$���k>W�V���z@�`����M�}d���eo|�v$�v�E|�SAo��1-c>'����g�d�����l�r�y@U�[���|�3͉��F�|u׃*���%�W�Y�_}[Rf�p-�� J$Q��Œؓ{E�p8�9�U4=w8V-2�R�x�e�%gA��?�� D)�7I5tUS,�P�M� +�P)H9O���TZuGB��#a�C2��w��ᅷ������6��G��h�e��c���<aF+%`�Һ�\f� ��à���|�=���U� ���Y�lF���Qc[��嘼bJ^�i̟��n����Z�y��o�]2ի/-JS�ו�e�Nj#c�9�xZU�9i�S��t��P�S,ovx���l��ߪ§_"*?f���''�̧�˫���l��*�2'�vi�y��7=���(�E�_��Bj 08Ņ��1���Q�[C�Z�baLCxR�a�mk�5��U�=X���D�����H�>��1m0�m���zF��s��ʱ8k]�_X�����/�A%�<��ߖ�
8���R�7ˊ���!�ì����x~!ާ����r��8c[y�;�f������V�4J8Q�I������{_1�|@�e��#����㕃>D�(�f��S����V���Q0��&�0��W�,Q��W������V�b"���77t�L�`5g�h�Ǒ�����uG�'�����H2�������y�x�AY��j"*0�5�n{�,1T��3�1n��F6iǆ�؉-b���Y�cL��>�������z����LfG��>?��p�_-�֐�m�����������q�z�2邪�� �w�嚽��İ�p2�Wdb���\�í5����{ ����\�1j(X�B�c�\v��⍎K��|��S@��n��iE>�}"y��%N���d~�(�7:�c��?[�b�L�\_��)�#s��袞�i��I]���' �NZ/����n�WHH��V�Q-mDF���P�4HA� P x@�KM?��������{�$�((>�(r����D�sd��IKw�yնbNk��!��'kc�/+B�X�Gb�=�_��Z�]�W�
��,���IC�QG�Dl�~�����!�Lt�,?+�}���?�+W�)��)����]��IGn��EJV!��8���Oy��TP"��ّ��)	�Ek�{�QP}Xk���n�`�d)r���S� �H���P,0���
�	�YSSi��͓2K�I�W�%]<p|DƗ��vѻ"��- o�u����66J���d�U�}��|�i�0b(�
9����Oe �c�������8!9��'?d�[ٽzᬩk��jR�x�
��l�Sj�sl�j��z9 �`qcӗTw�=��/A��o��vg}&�ɚ��\7���g�K�	�vf�M7�?wCSu��/��**{(ݷ~/�[� ���m0��*Z�7-�&�+��v����9�4��ό�����U�'�
�H�0|��y���^�A�� ��C��zv�����q&�?e)#�1�Lul,\��m��H?V3�ՑU��l ��0���
z/5���0�b��k�����O���>���Y��Y�k�.lbwB?ex�j]|r�3���������>쌨�GH�c�eu�h�xl�`�gM)�%�۰�L�6۾'E�B����5XVs����d���'���&'~0�R�r��\���H�[���t�_�g;x��K4�(�]{��w^W���f�A�?�{tJ4:���^�������o�M���k㠖�)�s�;��x���U���,K�ƻ@r{nxy̓4��TW�n��1�d |���Y< n��_w��+x����ζ4��9h
��#��x�h��X�~l^:�Ԃ6d;��ܐ�!��'���D�˾�4yR�2�wwZA��!X
p@*�<m��hX�tZ'�j�>��K���.q��|�t�6a���#fi�5�N�U��X��a�N�T�"o��A1��[X1��)�`i�Z�p��^{J4NG�l�Nn�@ϼ2T� b�<�V_��d__gK	�I��"�!��aÂ�p�Jf�6|^M�D���������h~�x���!?������}_́\��׮�&&�hkx6���+���5������,�<�����^#�寖�����Gl�e�Z*��h��mQ�J�?����!=����Cŷ��T�����.�����"A%*�tB3��/W��qD��Z(��߉�9�C��H%;�sa0)��Z�M���*E�(�Z��bS�L����&���kc�����c=�1���yJJF���P��@�,���X}����ǎ����y�G�!��*�sLj�I���|-��FU�)�Z-�P�����b��O�raBQ�Ln����\Ĥ����R�����c�t�?��z�E���Bͻ�p��=w_)o��������0'Ј�h�"p�[*l~��rՆ���󘒓�S�����d�[��o�/���$�(u7d�p�����J;H�,ى�o%�n�F.��yP��1��� 8 �sA�c��O����1����Yz5g;����\�-Q�i�rA�@��n��ַ=Ќ���bӂ���%�wN4R��I-�Tih��ZO�5�Z� P9�V@S������� 2�G3�t��8j���SѴ�2����}�!��_(�Ш �J
�>^�'��B�:��&����^�f�P�S�rX�v�F;�%�uP��)_ͽ\�$?f��S�8��u��i�
cfA�Fme:!�1��:sI��KOi"��@%г��:���tr�֜vS~|\��t��Ǌ�>o�Ow���r��)i�F-�!f�{����<�˜��[*�o� 0����YEL���{$��vyg+��p9�oԇ���_�1:T������7�s<�&.g0A�k�п+9���=�P.���|�\l8�Н�����IG�,b�B�|?�H] �@���*5��N�<-�"�
4���Z�j�L6y�
����Ğaw᪜���0�5��TY�����/m�1pB��jj-*�&%P���֯�Ę����Ds!�R#,p��F}vr��3�V��
�?m��.`�=A���U�6!�d�78 ������i���y�΁jn��
��c5�	��:�Uq�`�N�0�f'�l�L ��[�u��z_��(����z����?v��(�g�4΁q5��!�ѭ��X)ďU}��%��>N������f�fØ���	�ѷ�%6&��}�g���{�C�"n�6Fχ��h�&s\�x������>����">l]pD꣌~Ę=��=����((�N�x�\֒)GXZ�z�n�����A~���ܖ�/�u�q�0�Kd�-�s�<:�����i � B��-����(4�- TŔ�'[Sh6hsR���T���@ܓ6��Sd�q��\>K�	Il9>PR�p2�d��Q����"�Z2�;�A�+� �Y�d'YL������f(&ky�_q"8\'�+�^��13�/$�ɀk	����A¦����jt������Mw]�k�D��*I�;��g��v���Ƕ��#g�UlZP-b4]P��n�J�շ�6�%u�3�+�1�fP�`6G�2T���m=]O�� ,�ߔ:-R� 'y�o�L^oJm�+��Z�'��(�#$yԐPX[I)3O�;�.�D�
��ޖ�c���<��!f�o{�6��±;C��L����bz����,��,�n��Ǩ�*K�l��gH��a�Ц��&��j��-J�>�ĉⅼ|��kTX�ݨ���T���h�&�|V��l���V���2?���-D�������0�O��ր:����>g0q��D �Z4T��Dr?���ۑ�N���8��u�=��T�n �\�������UT��Y�2� 	ye�̼/�dj/�z�L̎��[qJ}M�����^��4F���#�:j�13#���X�'���t!�_�B�dW��4�h�q��Y"���a��=��8u��v��u�-���B��t�����r�.Wƈa�_�S��z33�k���Y�ۭ%�i��}9�]�^��F��7I�=b21ނ��͑��\�Y34q3Ya�{�X6a/o*v8�n�
*v��S�60F�z��/�9٬��-<���t�]�Ս�įv���n@�^(�V��47����>ޜ��D ����}J���)�S�Q��$��#s�XXh���P��*��x>e�G:�:dE%҂���y-'D$ٻLx�d�H���R�-C���"�OA��1�}<�����)�
|,i�J�㜗�bq&�ϒL�s�b<T �unO���o�a��Y^�qNZq�}�wcc��
��*S@��y�'�ۇ6�T�	����?�n��E����Ӏ�Ƶ�"ǫ�{��vPH6�*��Pbb�{���e��gW�:�A���8�C>H7������g�Ā�0:��K��-ZoG��ĥr$�H�����:0ӈ��{�]$�v!l�RlSь�<��9�*����j����`˭9�b���S�;�J�������4��ߵ���|�.|5$%>�m>�]��j<�yv@ztt,3z◚1C�&Tђ�]�������4v|�x�8�1X����Yv�\�{M�@�n't����F�>JB�x��2���i�鋐.�A	�ʯ>���y���v�@��b������(�#	j�����fTTw գ��M��ӎ %x�U�q�Lz��Y$'��$�ɝ��f� �T�ݜV&���z:��J��&gr22[��OP�y���~���̼V�����2�@�i��b�G��8������GṚ)�&sU�6no���K���"m��\��1���B6Yݖ�������҂�fK�����^�_Xz���7�t��%/�����gw��҈�S�Ͷ�����u�L�Lc��f�>B�i�`�3�� Z�����:�˧���zo7� 
!�
鑸~����_3�<e��t�������.'�sw���&S+��w}�k�8�9��N��cUԅ���h�����ň��p�����N��w�s�{zS����/��B4��j�!5<3c}�D[����,�dR��~9��{��Q�ݱKM���uр�L�h�V��dw!���?_B�����F����+���T��g=�f��Ie"@)bm
�Qb�?�ʥ�ߊ�<�#Yf�s1�]Fc�@KA0�:1�h��+�ۃ��4V��ա�"u��s��Z@0���v {�q�B7^z��<Q>�=�q��#F�sc�f���X�p6.��9~ �v֒ZB���T�K����p� Q�Zt�ۧ|F��˥�Z�"��v�#����R�x,pj[���P8=<�1�?/eQB,���&a�3O��ݻ�m��fd�:����[6㘍�/�t��]&��Jw��s_%���	!y7:&�G&�lˮ-Hj265x��p��At�>�
��k]�Jr6��
e� ����_��|C@q'��ñ-҉&d��lS�t-!5�U�H��b���j�A������dY���?�z�{�JO�3?�c��y�V%�f��?w�B,�spg���h'�Xı�����ƣ�ϲ<� �6՟����
͑�F��@��J�
���74�����F���Sm�؈'i[+��D̩��>}՝����^0F���n�\�I��Q��8���ڔ�>�J
3u>��BxWd�bV(�x����7���hUע�������m�ÓM�$��`�n��J7��h���e�Z��ݔj`v������w%r6�4O!�;G&R��01W0y_�a�?Ͼ��\�[צ�a�+���O�H4�2ѧ{ �	|L;;�����+|Һ�PN�\%�x�1g�p�:�1�A��R�@�?Y�~���B.�:gW�Y��Y�%�v���2_h�`��U����%��9t�KE%��1�|9<�8�|.D��GJ���ۦ#��:[�,{���yG9<3X�L��tZEԞ�4��,&m��Zs�;Dx7��W�{�qj���U�+]���IrgV�F���6d�Z�G�L��n1���Є���9Z�6m�
V���U�qRh�W������H�s~ux���7P���1������.7(����Ѧ>���ޝ��0�to�o�֛0w��J<;O&O�~���~[�8NLp�{���u��ls���ߏ�. _e3?�C8�~�6���Z�F
S�aVo�,(�-�蠷![�_Z�2�y��@��گYhq��j��C
	~'�<}3������ؗ�m�����X̟~�v	����2�zP#�y��J�-�Ҟ��Bu�Hv�ӹ�yJ78�j��5���U!N-�P��7sd�Q�"h�!<� �=�AB��. �}<��%�B����f���kz����0���7TQ�a_z�D��P-�*֦H��q]��8�H����|�)�`���2��N��-:���P�1^��a]�XxHe��޸��!�������o�K���m�H!7.sG��S�oz��l����C
$k��1�'�+����톲��=��k��;[�+���Ξ�^�s��.�$=^�-�dL�s�״b�N�%�AS��P����hn�E�q�vp3ȴRl�]5
׺\�R��ˬ���!컳'u����!��b؂d��o���qmF�z;��l������ǲ�������'#�m���R��M�����=�|��T��}"�ig����P���f�l�)jy-�3֐��w���I]���"�ov<��mU+u7xE%�z�t��m���d�;�J�O=� �@���9��P(T�+ޤ�/�	��H�e�s$�N.�D0l�Y~ޢ����v�{)Lv�s���^%�
Tn��R��90����ςw_Ǜ�k$R���1n^�������9\�C����p:O�qT��pwM�/��RQ��2>�i7}#���!��I�2��r��2�Π�4t�y)(�:�G��$ͭ�"d�̢t
 ��xj����x�uv�F[sh}���<�{q�si�Gȡ��U-Ζ�X��EP�_�gw�6�Rp��"�Q�![<8��
�������%�muz9�c�s� �,4�*��Gl����{�2�.�}�[��^x��ٸ���g��0����h��g6j�<a},��))��R��\�Uo��4�y�3�	�.�*��-=��CVIJ4��#����L]~NGN|2RI�6�_G�_n_�O��ni�����(�֘�b��%?�_4��E��kɨ
&-i��3�=v�eح���%�i��4ƫ0zٟ|W�Җ|c���o3�=�fm�t-G�)݂��p�h�kY���D�{�]'�8�8>����zSǫ�B�z�^?/Vqj��YCE�q<D���[��s����8���Y��hw4E����O�KrĒ�Pm���
����N1�	��-��_r�e��yY�Q�T��A�V�S�m庴��}*D��>��J�-j[���c��_jЇ�~g��Z��\.Y�̼������b��O,��P���o����|vL�с�R�"��$,DQ�-�,�D����%�����!��S��0�;����:F��,;�*oA�6瀴O�Uʢ$�(�ƌ�a�9�;�9�m�:�{؎�>����P~��oD�Z��g�+"zX49�>98����D!�S:.�~��У���]�Sq.c"ϝL�]G�N%���f꠫�f�qZ@N}2����"Y<����Ԫ�%7��
t�?Bx�|��BAV��	��}�U��h�Re��%�� �����|�@	�-����լ�w!I�8鄤i|+�i\v���M@��B�����9n�¿�M��o�ۆ&{P����43�·�	�Xų��V���*Gp@���ⵄ}B��2`�jA2��9��	>��U��W��!V^�Me��3�@�/J�P|��7q0#nɫL2�?Ƙ^��qu�>mr��=����_�dδw!���$�9T�&�^,'@R���٣>�M`gW�	�đg��\oy�]KZ����;f_���ғ#6����st�f��A�$pӇ
3��L[3���PΎĺ�zCYo�Pi��F%�$�w]sȩ3p�{%V��eXW�IaA�rf"���Ү������ф���/���TI$�����݁��,�]���]��=!"�Ѫ��{6�!���{��� �7�{��9���my�_�-�����p���+鬯�獗��z�%b�?T�QDr\�b��1{�]���������WyCp����t�i�"�c�M^(�g0�M�5����&J�RՀ�6j�dBe�:�@�zu�
�����#7\�	Z�u8J�}��}�I�G��_��yƲ��#>�F����S{����b=寜�i�I����\,��ˌ��/�o�6�PU����{�䘰�6�mq�p��2�'��4��b2 V���{�����w%>ݔ���uX�0�YR/���@Z�Z���n�K3L~�}\�y��/(Hj:�K������'Vtҍѡ��vWZ԰�8�a�R�C�̬��]*��,z���0�M����!�Q8�'�|��=�%#!^"�m�#V�Lqf�y[��	�����eb<Z:h�9�:�p��V�"�Xɵ��1��I>����O����N���T��5��/r��?���)�>Dy�[Y'��@9+�3^���cqݤ)��1��+B.� �Y2Y���r����dz��aݼ�(�s����B�/�GBƎS�î	�@l��i�TIC�˸|�T��E %���2���Pn�`�/~�ڱ�?
�2JM�ڟ��n>/�XH��Z���3�q����K��g�|#��*;��7�I��Yt�{b��R�W3St�u��QL���Vs^@O���p��Ɠ�����Aw�y��C�X�����͹]L�����.��ꊣ%B^��FU&��ؒ�1L�>�췉��P�ͭ͹-R)<�\���Ҽ#���z$��$����U�ݳ�o�3`TZJ~�o���WES�����1+`��/�;��-��X�oO����6��ԟ���^7%���=|?��(�γ�<}�H�S0s�F@np��h(c���.���S�$��D�1�o7�����zU=������� ������Q}ϰ[#�/y�:1B~f(�͞g��[#�շRYP�W)�d�b��c(�[�:)I�L��%F�ǡk� o��G�[���'l�
��2�E�y��
���<�������%dŮۮ}#�S�f�_����wFK.��c��L}��gc����`e�+�d����2�I�N:��d���U2(˞�m8@�R��=�7�@� -Ɖ���u�Y�M���.rR�y&�F"�ܛߙ�T�2�2([�>4�Q��!��+m4��s�����ל@E��iq����V�xlIy~��)>�R<��6����!l'83L�>���8���䛭"NXu o0�q���lj�a������}�R����ˌ�*z�m�c{RJXk	=:�)�
iB�1���~��Z�t���FS�ONxЃ>�FUj�*��/F�;%�{� ��-�-��;�4�����������O��1<���+�TAiL�)�rg�ŷ�ZLy;
�#+}��ok�
L �Y�0-����΄Ŏ���6���{�b�bd�<^�w�3�+dt���1��[�q 8=��B9o%?E	�>O�~��|�#+$�ެⱩ� �Q��1&�#�ߟrQ�4�=!����>s_��²a)�� �x=��q�j���yH�8y�3���o��H�j�^\�V�M:�=X;�m.)��
��U�!����x�޼)	<뮃*��	jK�^d��:=7D�-�b������L����&B��c���Ќ�<&�����4��e�#��1=S�:2�%	p���@b�����b�\��Сd��U���p�P�Q*.$P_VD�
�Y~S�5�$hP�&���Z�\y�G��Hr����ͧX�.=��xH�_�-ӫ419�rп��R)�2��{�fD-�D�յI���SN;p��y��b��r?Z�[�T%���;��]4�w���@Y���?��Urj��Eߺ�w�O3��9��k��J��8>[��^���wGQ��wn
��鱑� ��13�P������^�9�EĊ:ĕ�D�]�o����;��:��t���+��?'�2���<B�� qp�I�	��*pڼ�]�4R|�������ѻ��l����wC �tEڅ@y�o޷���ٿS�G{���d����w������W'D�Z�� C����s�4(�ƣZ���Vk�D�'�:�E�g*wuU���y%���d(+�-�_�����	�F2��Z����ʣH�o8���MÈ]^ʦPs�p�g���QE�A�!�#���5(�����m����T%�Ś�9W%E$�%� ��9D
���=�9b����D�D)���̦�x��K� ��q�U�.��N�qRTc	U�u\3ȃ�o�6&�	1��H.M�}��P��M�A��G����CHU'�������!h�5Qj��O���Z��֪4HE:�-�`���*���
M��O�kA��I�pS��fB�P����WS������I2J�#�?��	��h�Mr�:v��-�}� t����-����e�a�8�4��Ͷ�o�N�$q'��	8���k����ǥ�:
������.N�sif$��W��SC�9qC+�ҕ�e��G[�����cw.��c���C��c%�PmČ�]y�%o�z�UJ͚�`r��wc��H���V��9w�$��k���|�L��;oj$l'*�ag�v�9Lu4������ �?��5���/���f[���F���~��I�H<�.���&�k�[WgI1ؠ���H���jA�xd4z�u$&t��t���E�L��H�LK.�9	yT���P�� -+���Ҩƫ!�u�V��X#��]�����݆�,H�e�p�b��e���6��s�K��S`�&)�7�Q= ��47�QT��Ԋ�G� <E�`,�z��Ć���`�J�=}�m�w��f� VQM���Gk'gV��3�O�M2�0n���!��n��៪C�4E�M�b{/��6�Biz�ptb��@�r��zZ(_S�{��uK�B�!m��t���Σ�ȦV���]˹z�Ħ�/�ad��Č�:yb�)f�YMeN^�1�b{U�8T��$k<3$�GP��`���H9q<��7�;���7ń+�O� #��GП��|���J�<�Rxb��¡yh
fY$ǧ�����aO���Q��nb���(�V7�҅�e �Lz��E���g'p������r�y��q�����C��]d�#!�\-��Ƭ������F�h�!�|Ժ��u��~.��X�-��J"�ұS���dQ<��k?��jj�hm���<����_4n��6h$�`Rx�jD�Q��5:8/���ϖU�Y�Sh8�s0#��cv�,*���{��"�9�k�0}:�=� �b��_Ԧř,_\f�t>�� !�:w��'�7q������e�A����!n�"���
�C-��6L � >�_oF���h"X��/�y�M?���qv�fz���m��������9^G5Q��^�A4(��uLU�:WRiD����/��<��L�!b`m��S��eZ0y�s����0����0uV��
dk6�evүt�s�|}o,�0�D��/�f%>0��"�/O�@�jm�s�KE|��Um��B9�����q '�y`��8Ԫ���\4U��L���O �	4{-�u��3��j3=�QF�=�53e�es�	����A�ΎWg o���r�Y��3��G����f�#x�:��[��a����&�S^��,ү�JhL�>2R�G���v�D/�
x�5Qb�����lϺ(�V��ۖ���-�����}��T#D�U���	Il�+]EBF��Z-V�S9:%�Xױ8eb@�T����gVe�Ck�/{�|�$���1�疻O�B\�KH�3ōV�l���9�1tLF9����c�!������0sX W�����15�� �'ؓm����釣�Ӟ�;__k�v�����_s���s���eř�v�I�,�n�ف�-�L��E�,	�����h�p�z�a�!�+�S��A��� �c2���'�0���w��u/�*D]Gn�J� ��ZpJ�Lhٱ���n���ӭ�Q'97v�S<y��֌�Uš&"��F�|ݗ�|D�s(z��].P3�&�f!x���}�M)�M��8�s׷��Dc~�$+���g �"6RIܒGJ<^��!7�s�}POn˪1��&�Ɣ�Rry�]�A�X�����k��(����H��
�LE��7N�����W��eʻS�Q��)�Ѣ�&�%8Ɖ�����h�qoB)sKWa�1X͙^K3�f��\GS&�6Pʿ3�~��U�L�7;�^-����Fy?l�X��l�2HuE�\Jۣ�>�C.����l��ID�-� ��4�7�4n|�'[�y9A���hb�s�#*���(%$ ���c�X ��-��6n�e�=g����/�ZcIֶ���)b���~i���o�>f���Bѡ;2L��+^}@���Z�U��,�{��T;�?+ni�'Ԍ{��$'���MXڨDG[�.���V��a�;�)]"s�͈Nf��,��_�굿D?�s�	9��y�&'�6�&</5z��ߏ��b�~֝���
�9�]2Ӥ��P4G��R+���W���~�1
m4c��7�*��-�Qe��!q6�a�Tݘ�0�ܚ ��Uz8���_��9��U�î�S�����<��zy��cIb>N����{
�}|u�MA�޼�	��D-CJͱT�:�ٍ�%�玑q���$�{څ�sSꆎ=��u���v>|�*�h	B�D��'�*�?�]	hcv�w���=KD-��!������F������dz���\Z�)�@8���ʤ�a���DH���ϑ|2�����RK3�><06��o Ojύ�'6�U��D��^��A(f���C�m?��H�"�x;7���6�f�~� LŚWj���sM�30�����>���[.^.��ϡV�/�!�?,�+f�����|Ar_M��(/n?��f�GJ��)��Пd���<���r���ݷ�Y��F�Lz��r.
��]��˙�1����3Ԡ�1������ȍ������%-,(J�l��0�qM�"����EC�I��@�k�7�>V%Xr�.���x6���^���B�^�)1�<��q�z�޾"�|���Hd'B�~����@�l�rt�V��4^`��!v
��P.��[12໠�X�c�����q���������7���ޓ�B/9�tؗ�l�l�_�s��� �X��f/ؒ�&�ꮝA�
:�f袣�4u|�H+�	�sٺ��E��=��窉0kd���-ũ�)�<�����thD
Gs!`�U�i6|R�y��w�4=YR�#l*�Йh1Ț�X�?����.g�ܡN)��܄�DtN/M��3���J��p���^hdR�z��Sا+{�k�vB	�2�p%z����@i��q�E�#w�*k��TC.��h��E׈C�1 �z:=�������Y[M����o���FG�5��y~�����Z��W�ܪi���h�1~̲�l�}P^v��������'6��s���B��q��<�vHfH8/!�9K�?��}���J.���Z�E�����J�K��]����X�o~oj���e���I�Pj�6^�y��l�%��}D�}���uK	ڴ�-��E�nc��憽K��k]/q�d��4aˆv;K&_/���U�1 �����ȃ���!�9[`�8?����݌b���Tw�PI���G��[��PWS���`��8�s�{�bp��3�)��uW;��4f�.�O�$L�vwL���N��
�3TŸ�TG �կ�Z�!��_�Ⱦ	�)�i� f!WD�>z~g�m��%��<�^�̜{�. =$��#���=e�Jjzx�9Ib��ǟ��­� ��O޹��H|���N�$?�5��Z%*o嶐/��6-NX3��F�7�U+lr�M>.�X�Su-�J�''�҈ah,�Z8�Z��Q"],S!���펙7A6��aX2v����;	��h�F�E��?͐�һ�jJ-��!x��	߁5?�MM�Z�㧛x�|C�l��I���h�>0�QL�ж�@ ��>�?��J� ^/�ͮ��S�a�Ybe�n,2;��%�DӶ��H��>��/�ݙ|9�9�/'�<|�>��ڱ��s��k)5'�� -�9����RyXQ�N� O3V�ϥ?��_͍o���<Oxǚ�<T���Ŧ�o���3F�*���%U�&&�p���`Ӯ��J6�ە�8�멏*ѹ��p�FO��07H�3":�`���^0�u���JUx�T; �}(-�F��-)!�pY ��ز�� ��9N�~��tF�� "� ��_�T;Qr�=S��iG4~�l��|���_�G,CzB�d=�����R�֏�Ts҅���k�N9#�j��h ��/^Z��q��b�^�-
*�2gli���.ot��O�J�\b�)�����d�nc"|���9�\m���D������.D�4$&)��!�RU'|�i�=T,~��'4��x��a��b�L��p�dH:��P��)�o/�"I��o���T��&���b�C�Yԥ����'�8�fI�@�x�:�����m����ݟ4���fe�]uYдs�%Ri�)*��MFk�>.n����[���Ս�.b�v�2=ff?B�t��Z�OO>�-�5j���h��\��'� ��}�:��sc��O��΋���@G����&�ȃ��y/����ۓ�POV���݊�DCl��eKT��ts�|�:ֿl�v7=?�Ď��9��(�u����C[��͇��~%���i%���0@b�sm�u�Sh���K�.�i��Y��$Y� r����%~軍X�rp,��tA�7�#l�h����_e�-�p����S�wp��	�`L<b��٩9�n`��!
�
U����!��2�~����|=59����W��s�8b�}��z�y�3àߩ3]=)��f��/�3v�A%&So"c�U�Dw�8{É�i�4$�YNZ�<���O�#�hj�ir�yg����!B�3/�ow��r�ٲ��������t@�>o��;�he�ֆ��Z�ͥ������O�8юN'�j�1�B�y�/�{�n�^���3�N��R	�1�������;ufݕ�����y����iM�`a����i`-�� ���J�2@�y��{djb7��@��q��Hm����p;�!	Ϭ�<l���j��Y�*�\*E�PQ�R��/�'�W\����m1<U&7�!@�X�-���'�狄~g��� ?K�iy�w�sZh@�w�����"d�v�r�~��J���N=]��*jW?��?�0�K���+9D=*��y~�u��kTފ�z���
']�l�NL]b�5J��G���)߬Ĉ�{�΃�/�ڥ�p�&�����v��k9����k����E��PA�Q���潔CU��,%�w�ecSվ�K"�ճ8����������'���;�djՕ�(�}�s�r�v��K�'6��^�qʩ'�L
�@N�+�6Ĉ�^z�J%��$X=�˗�y�i��&�'^��>u5�W�N-^R��R�ERD���#��a��0��@v��n�K�*��W��hN��.��:��B?.�O�j�Z�0�(�z!5���Imx~i q��|�
[�O�*#r�>�?qwG� H���L�L�?�,w1��J��P��T�?�q�'<.mX�	渆�?5>r�f�q����R|04W}'ysC谑fÍ��8*G龂�r �=ݘ������8 ��g_��`�޺�
w6[0��j�a��aJ��7�*��K����G,��qH5浄�+��Try�އ1����j����p'�ݼo�OL�X� ^��$M�s��X,��BYu�<@zN43VZ�� MthsT?���r���We���fI�/��'���ȥl�H3Cc�1�2�ݛS�Ӭ��
��Jڹ�t�VpS��w2�#�����+��7�ը���dJ��W7�?4&ΰ+l>�$�`���|$�P�k�+�Z(n���
�L��)�8�A����� �"1�9���fh���D��tl��sÞ�?u
�b�t���r[�k�ܞ6D�Z0�VA���,��G]YO�q2���6!�W��m�\`����Q�S^U�rW�Y��̷���}��J׍�S��I�`,��v�����|���1�A��ӂ-8 6�+Z��@4;���aWa��o#���.�19���W(���!k�u��R����t0�=�.�ϐ�Ӻ�y����-b���a}_Vz�����L�����)b�g]Y��$�I ��d$��3�e���d�	�����>��^給֔��䔂R�*X�DŎ��� A���s�?�.�f�c�Kr �Cd��ѷ��6�t8e��a�qI��(�J.����;SMoB�s먻*~6=�`��xW�Ȏ�rz�C��3�)A C`���c��w�٘A���l���2������W|6b���ML)tTU�4~�~��2����7�����T���8�isX���D����P6�H#ó�̓�CR.�LPR#w����a�f�@�L"�Lש�h���"��3�6��_vy����5�� ����/KaӖh����ٕ��6LZw��1@B���;�Ǣ�(/��/}�u$o#�b�=Ӄ{]I%��H*�u���ˉ�_0t�w�P��R�^ݚC<.��ɶd�o�U.ǉ\Rx�͂�t@��D�!L5;��䀺,��Z