��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@��D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6'��4��f�;�J�鰷:�ذ����?�R������Ԑ�r��ZJ��1�8c�č7n��MQ���������1������CZ���E���^��<�8��7����T.�nO0$�MP������m��ݪ��2��k`0nՁBD��bYWo�2C����v~/����P\��N�Ȭ��,R���rHx����b.�z��x��˴�C�ya*�gmӼ��q�L��>�Zb#\�R���|��M�_���W��9��2v�uv�R��q_�Hz�~�����XT���AE�`�A_l���$A��y?!z��=
W��&<]`B�k(ՐC���5�g��9�8ѲRטY���n&{�F"�[��ChT2FI��uWo��.�g�nҿ)�+P�1���M�������P��O����p�o�w�&�1e�>
�F�`�۞y/*�V�mj�d=���ѫu}]��;����Wz%ic���h�ڛq��PJ�ԟ%oQ�ٹxW~�n���`�E��2���w�����������wD���^z�g��f6�!r�sr�]��w�'�gI��	���ܤah��Q؞U��������UA~�b��!֡�a}�O]q��-�J���ڰH�w�(<a/ܠ\����U ~<G�Ԟl�N�����SWi $�!�o��	8+�p�� 0�N�d:>6$ zD�i�Y^GxD��<�L���P�tÔK�]�h�E�T��K�Y�r쪓����_�����^5-oڇƥ
`fOd�ui��L����_vS�k�B�����Q��w�v��|@�p�4P�f�����]FV��;6i���a$F%�'_Yx�Viz=�/�)C6���U/�PT������m��5�[B����"W70�{�#��g�T��nF�6�w��H.F�\�P��]�j]�4a� �_�i@с�o�fM��3�����<32.Q�?X3��\?�%������q���8�Ы�j{�=���o�/��2��b����OV�<mP�OV��Q~��fD �YmNiT�)y�֘����q��l���9�n3�D{G����Ai�U�����w�}!RV���q�I���?Q�"�$;I�i��o��j���c(�ǒXΟ?K{���a5�Ws~�`&�=��Q��z& �cQ��d�Cw3�`�F[�:��`m���V��6��v��@�f*i�с�%yA�m%⣽�.�*�T����e+L�x�����a�ͤbMEFD��{��#
Z���mQ�xf�z�_��my��� ��Ѭe��eS�$-i-�&`{�X��Y`�s����t��UK����w�i��G��)�W���u����U���6h�b���Kp��PP4wC�V��#������ֺ��{��e���&��b�3/�:wV�nf�h�����kU�d��{�ny�_BW)�3\��R�aa��aݳ��c1���l���8o+�N����Z��3�	z�Wʗ��/��&xA���:^Fǹ����~��^�W,.n��(�C�o,T|�h�S�M���"={#�y����{Q����Y��[	���u�@[�y�0e��c�w����V*��s�F}K������{}�;�	o�1ƿ����G��z������Ny���:���b�3x;1,��"��`�Y@�v��o�φ�g$N�cp!
�f�ڤ���~ɤ��e�OȞ�Ȅڷ"��Np���"ȡ�
����T[˒D�ZL7�!ȫðԪ\���2h)
����ʭ�O+dhN[*s"����]��?�����W���EP4�[��U0�̈́p|=8Vǘ`J�ij�vV`��ذm%I�֛�f<��H�A_"�A=�Q4�T����H�~f*Zt5Rlҳ���B$ ����hџߩ�K�Y�K��C�OF��Op��;fPeUw��U���>�
��O���� J�?�eL��f�)�D�8�&T�0&*�߽�+�6���{U��1�r�C/pt�#r|r;��M!���^�Z0aZ��K��i�P>*r�_���͊�/��c�\:@�P^�b�Nd{�P��	2k��4|��R�h��S?v�-p��?k�z��!lB��@���B��@��9Ӂ�C���F��]��6�۝.{�M��d9��H�X�CO@�-ו�<��DݓD�>׭~I��D"���s����WKR4k�y����&�ߵ}L�ɬ0�s������Vv��p-N��"3*el�7�.Ͷ������ON�R�kTl�H����.#g��à��@qH`��X�_۵@ ��䦁U�/�	�ݻ��!q� |R�FK[nܢ��h��?��W����|�"��� ��{�([�w�`;[��SL'���r��ժ��X��p]����xI��� l��յ� � o�!$�b���lg�%�ժ@��)%A��|�5�C2%Q!y�u�2�7���t�wG�>�V�m�$���|E[7{I��x�l�F����1��<����+�o��~�vg�(����uT	�c�I\����1�4�r�0t�Xt����_� ;slyd��7�Y?#u�=��ay��;zo;F8gL#F7��o]�gA�g��:Kǒ�ҏ�Nc�������`�WY�����-���֘Z'�o"����
�M�h� �P���?��r�"�~TJ��n��(�@'�TJ��r2��I���vq�Qk�4?�������7ݒseFq�����6�&�w��1�����'����*��V'#A)�^��CAX`�y��.SN����խK��/flW��iu8�%9@X}�H��A���zJ��OwB��K��ӈ��H4���l�������͝sP1YQQ5�a���3g��9����|IoˡT�3�7q7�hx��Kp���ua�[GC�ԃ�%v5�����ɋV�X�~"?9��;�(�"��u�#FA�fC���ķ�B��cW��al�=����V,汯��*�z��u�j 6To�~테p\���z�D&Jc����H�jc5Dg�p���.�a��%>��^z��6u�0$�|s}�uıM��PKB��+�X_E*AU��i��j���T/��.�C[���ǔ��N�@j爽cO��&B��n[N�f�.����a:��6C0�����F;�dLo�'���#��<1��������GF��N#ͬ���s��Eew�Y�-�S�o$p��װ%��$���j&1��#ӳmp^����͜�����a�D�5/���H� ���Ni)䰫'#�Dm���r�
-�[�Ƿ���9��g{�x�Z����cdFRe�S���2.�����xB�C�V}}>O��+��׽}�6��w���v(,變N_���� �&֎1�&I˦�]'��$	��D:�_^8m�X����R�>$,�QX7]���ڨ9�`<�C`C@Jh[�,�<Z�W� QK�f�8�����_p+��su0v���y�e���bV�z��m���@�.�r��jy��Ǚ^ʦ��|�|��5�� �ˈ�`g$fZ�����h����hqJ�*@��3x��c@h/|��3���!��&�cA������uS�	w�?�Ks�s�d�!GW��/v^�ו�u	^*�/��C����F�
y�.��J�"*@�Z;U����c�l�]6l	�� �Sdp�m���j�9��BR��m-U2~��f7�˷9ȺJ�~��'��b��:N�n� �7=8�t��:�U�|�:�T:�HBx���n�n�L1R3i�\�Z3j�.nX�����X,�#k$�DVB}׭Ԯ��D��(��y.f�Х4庳��J�]L�9�,C��$j7���vx��9?	���?���^?ى���\�Ց����C,�1ݮ	+�Yy{m
4v���ۮZ���t�~Q�/)���EXD�QۉP���	�{/�?敔1��8m�>T��t�F���;���������L���������~p���ؓ 
FD��g��60BRjt؝D?�I��%h��">C赡��S�ŋ.2��!��c��/.��B���y�s��߷�2�:�A�ݩ�.[X���6��s@S+S\���E3e˃�b���׵*��<��z�tO��z_-M�>���k�����p.�9�B��5=Z%l������q�Z�H�w��p�Rœ#�g���������JFNG駡쌌�KaC��l�9ϡSiE��!������=G�~��>x�uÆ�r}���Z�_�f��Mὠ��5�(9��� k-��^�� �ɓ�f�qw��A�c!J]�O�?�[ǉX��������5���xB��萻4�H�:���X槗7�~��w�C�������%��~*�^w|��M�:��EU�--ZsD��PIng��I:�^�eX��|f���;�-:�aq��>�Ө�|�&]#*�:*CF����擏t�_:���KT)xf-T,7�W^��� v��I��;�O�E~��{���D=����-���Z�ʟ���y�rJ��3sn��D�n�MQ�1Z��ial��������Lm�bY�O���"�	�GY�����&"S5&��_��g�����k��$٢�2��Рԓ�v�"��Ѫ8�>�n�c�ǜM����w��b�.��`�vRT�3Q�Y��!AP:Hy�~	�/��3k=�KFa+Jh'P!`�f+X�u\�z�
�hgU凉t�{�D�E�e?d�~ۼEݱ��Q4!Njw�}ii�j�f�cXve�_s�U��g�rT{T*y�3VM]<�F�7nD �'ֶ=k�/%�V5�F���Z�E��k�ȬFǨ�h���d��,T{����8�Y!RAOL���e-�A��/@4�����n|Q#:dT�>9�5�'��,@����f�<�.8�V.�+��7n�tםӱ��R����Y;���Tzr���Còδ!���w�h�A!w���JK�s0�ǣl�1��W(��8/�*��}8#ME�d,Ԝd{:N����k��b/�E�j �w�_���C�`���"�^����"un��C��*��ӾN4���	��l����pdK��!��e��v�����輍!���������/��+���뤤��flO�uc�l?�Z!�:�-�������[���)��8��o�pd�뵗p#�.��MU��:�}�0c���$����BN!�l���aL���C���ُ��rA��}���kI6�/��Ŧ�g�E�9:o�m�ںU�2�7$�'�T��F�J$av�.ե�惠?�E�_Rf��<_;2/U�7�F5Z��+G�����=���@������cQ*�Zd'E�7,���n�1����'G
#�I��!�M��)V����Uy���!f��y"���e�q%$#�D�����!�b-6B�X��޷v�T3��=IWg�$����l�+���%{���z���1p|�^�	�����ؙM�_9�'k�8���qA�W��<̅�R:��'�D[��JF�Z�}�3��6�i�R���+,��m�۷�[d�ɂ^��'vs�֊�;bk��&xtw�U�KG�=9�k�!0K�ӹ8^	B;H �`lzf*�O����tm?�0vQ���@���g�L��_��(QSU�P����h�B)�<��<U�к;�'.��OL�:��L�]BS�� 
���rPԝO?��R�sJ���;
&K��YO�
�ч����CW�@E5��gaNQ�K1x��*�(ɆX�fS@�����ϡvԔX#L�ǅ'��-��w���1�MH\��>_鰾[=�x՛B.��Sf�8�O�|�Y�x��$�uSv� ��g�n�Z���Ţ�. �M<�N�Z���R�ĕ�?VVc#RG<���`�X������.�Y�1�O�5����6������N�p���0��A�P'No���-��f�g@�
1u��	"a��P5�f��
�OA�i3���0�k�
��I�ẫ��������(A��Γl�k��I��� $�e2�W:��bZq2���ԋ��\ ��Ҡ�����.���Yټ9F�rǕ�>�3�1��v-
to��Y�^xv֭��8�����,(?�)�"�.�uanI���7%����$��������V��؊��1Tx��j]2. \��`u�Ū~�r�]1Jv�f���Sڥiq{�N�&�D�Pz�!�,I�.��ͨo��ܾ�#�w���n���C;�N9R�E�r1�
P�U?�~p����&۴��zɋKw�� �jn<<��f���2���y}y:����%����	Y�z��P	Y��0�zho���h�����+T�����5B�-��ĝ&0�C�,�<��w��* R"P;)jO[�|��f;��U��<����9�R�`�	s)x���~f�z^w��T��?o�I���pޞ>����L��a������;G��d�
�莗�L��W*j�R�6��%0�
�Z���<`;� ���?��Z�ƶ�gJV}�9w	*}�׌�k-z�f�Ի.�H�����ԧ��`��9�4���w�~����F��β�������qIE%����(4k�[���8�	��Kqy4�V��i��jk��e\	��
x�C�#�=t,�i�ns��z�g�+���q�x�����v�dӶ"���)R����8B�v/J�fPd�,C�VN�{։���J�R�$p:*���Sg%�q���N|��~�����0��@���]K	�T��5�~�ӿ�K`�oC��n%?]��^az��!J�Q$������B�*ߋo�L��#0n1��f�)�4uW�˟�dmhzf-�����R�x�J�	��IX�����+p�����q�ס78l�2w~j�P�Y������n��	�N��~�����5J�8Q��&ȭ�`�g<�R�zJ)ΰZ���e���]k�%/��o�	YI*��q�����ϙ�#���,;m�δN�F
�t�E� x����7ՠ��N+��Đ;feO�\(_q�C�2��!8���~�b�~y`� �7�Db"[�!xa@s��VG;JQؖ�DX8^�x(F��C.�8u���6-P�O���h4���S, @ꠄ�{���@�!@�Z�*�0�75���
HH��.�MV��Y_#����7�R�3q���%�O����wp�mK���A�Q�6Q�_�倉N�O��E«� skп38��ID`-���N��k�F��y�$�:�G8b���ZϨ�p��t�$�{}�s)�#�!������u;�O�O��~#b��7r�PQ'�������!�I�Vd��}8��K,�%!��Cmm_�o򹷞�3��u�w��*�k�[����x�h�3���c�<O���0�r�Ă�:i��;�*��kJq�V:j!��3���Q��*H�$��K@�^��n|����;�������jxe!��ch��_4���f�l>������˷��Y�|���ǳ=J/b���VO(��8��\�՝,�+*�n_�a�w?�n(q��Ck���i�N`mv�Q�1�\m�(�C�S�^M�$�kr���C'+��2�$)r�L�� 0�Wz%����)M��ݱ9��.&���k\˕��m�P+�˒�yGH~��1b���x3$p�`���o^����X�W�P�߭O�3����p��c���"Z�MM�:*�m��+��3��6�c��ZG�7�g�"w�<Q�דx8Dd��u�+4��ܬ�����[����^E+s'��%��;3qey����7�ݹ��#/Yyla%,JqH�m/�P!|��Cu�}@h�Y(�Ƈ�Q>�x��$��k1�-������>v����"�	i&���qL�1/� G�Xg"�M�sL>�78�]}eϹ8	�ر��Il�dZܟ~�k}�mPQ�s�!��d%:�%�.�3ӜX(F� Фy"7+���eF�gd�w�?�-ܶA!�)]i�N S%���$�y��O���@7�܅���qo	�G�%�И\������W��}	dB���Z�-�H�m=�yh���;[��q�6�`<���CQT�ֆ��h�ރ��8�/�,�a@^�8Y�Y�l���10�d�R�g���Γ��f�=x�*2k���RƚL�F��B�KW�W�cȆ��|�d���8�͒_��1�7(V�1��b_��}{W*^M�r�iGaM0���b���|��B�'��Y��kI1����.���s�d�&K�2�)�B�HkϺPw���w%;���}TRQ�L3�>pf��t�����uUY����`E��"�@�M�u5��&�9e�E"����+�/���s0P� ��)xƧ$۠��։>]s��'�'5������1�_$M�R���w�C��J���h�x���c
&�Ď����P�2
1����@�Owo�=j �(�]G��0V����E2f�����/fƝTX������)P?�M�\-���Sf��a'��F��Y�'�����9cw�ӵ�˚�6��搃�� ��@�7|�����ױ�v��k��VkyO�~��lA�r���X�����?C�lI���l5$9v�c�R�P�FSt*)+p�W��f����13��ާ�/��\�}z��ݹ�wv�0"~]bO��S�	i�a>`l���A��.��n����bX۠m�,6��Xr#`vuR�K3�c��n�S׶�
)d���&PE�l�'N�f���g<���'>�gY4��>\�Fy$93���;�}_��  ��fŕ��tHL|G��ˡ�[��3}m�x���<���mc�Im��0���j�����}�2�M9�Bqo����
!p�6�X�f�ғ�ބ?j�Q�G/=��
�+~����"kV�\+��ǔj|�q(��s2Y�͘mг( �f\b@��/�����7���Q�In!��EE%F\�j���D�e'����ls��~+��&��������� o<T��޶��Ǟ'�ڜPs���U"x ��֦3�դ*S���Ch���x@�ͮ����
>f��كc}��I�C��8a`t����:f��F{���J+�7z��t��{]?�߲�[��$*z5����8�ޯ�VT�~�D����54�)e��Z�N�+���0�K���fJ�Pe['7$U�|��Jn��W��1����i<:�/ɧB�,�)N�f��<���?U�G�]Zޓ a{��~�p����)�r��G�)�+L<��ثO�3�"<d�|\R�8^�ߣW3�+��:m0�!��x�z��O�2��`��=���h���Mb�~�u��/��$3�gS�C�4z�s�����8a��8��q���L��{.�*�(��]����'D�E��n�T���@��4�������#Ia%pG�3��g9U�~0Q�>���hTh}���H��򎆚��k�'p���R��,ƃ�&��?�J" ��c�Kv�_��M��k�OȊ=Q�V��t������᝵}^��$�+**I���߹��-���%۝[N���M"��$��v%����q��*@:8�0�'����nbQ��f�m��0�ۺJ�U��$�mY��� �>W���B~����ߵ�Ef��� �q�`�A��Z+�|bME�ʱ��PuCS�T?RW�%M���ᙼ ��/j�n��t�������J��KےV*����j�Q�P䧙�R�OHf�#�vve�;N���������PDǪ~X��8�����kY*�H$���|Y�ֵ>�ކjns<"_wm󔭜��z��@�P$�*X����m�:�ˑ:=�ߑ���� Є��)_5�%�A�>����Z~w.٩�EZ����]�����}W7�3!u�Zy���
�\+n~����v���^Urr;�=������J(���8�#��q�����+B���TP������.�