
module DE2_115_SOPC (
	clk_clk,
	pio_led_external_connection_export,
	reset_reset_n,
	getmax_0_conduit_end_datainput);	

	input		clk_clk;
	output	[7:0]	pio_led_external_connection_export;
	input		reset_reset_n;
	input	[31:0]	getmax_0_conduit_end_datainput;
endmodule
