-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yrDRaFyTdGnW3NKAZckaI5yEPOxvkbCcdEnuTz8mj0akdHm/50r1U5fXhN8aWd84dVan6lJOWv9H
PpBgQQWGgPdt+Il56tQ2KCr/3nA4NvdFYEkdJ7MIZrd64thsJEVUEVqz/hx8L2zTqJo/RMzghXM7
QdWmj0G6ImZCDlJErw6IZwXn4FFDtjyOB2MP13samCCTFEvFCtWQL03tdpf4vbLGqJu6no4cOZpf
OsLGzSoSt3/UlH6+N8ODXLYGK6a/e2duP2I8++IC7Q53LBfaABhclMJJ+vPc0rntSQbPqDDp5jS8
GxPDHFAKPy3kB2UTZj+qqul6GdqZEQxgFB2AZg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
RfgmA7vttLI1krAr9d/tIvSQV03SCfdjW7/nhX6GdVBTSW//PFhM48xivezC/Tin2kTc3gC0R7s9
fQevg5eYAxkIYu3TPITXQuhmFwbMsJ1mmfnyxnxghrz+4TsL3kTmmLHcd0/jCjhc0wCRgvi6MCKQ
XVKPjoSbUvOf7herErlwIi02EKBBXmP2mvUH7szJkSZCvlQtfAM1ZmG8M1MATTS+2Unk/q5BXH7V
MMp/KmZx7gZbnI/ejzpFmR6n4NxOa4cIw9JWsa3c6u+zNGPagQhU6tkzgxj0fWqi4G/V3qwsU89s
e+epLytR2anT8znXWRQ6FGCNSDDpmRCgMOcuoUFNTS8KPbZjO1AqrOBnxzt+H3Bvih4/8gSuvPgj
GKsl0/pVyyO4peI4TX2mT//vZrrAidz/cptuK1ruvz1lqfcQZ/6Q76uWtvonm9Lh9xdTssk17pJ1
SuXhJLNtpVBp9yjqSiE0DOuhyRwgfcVmPpAPqzF0RsjMgi4eAgZU/I9nF/kWVXfUJGyGSp0M75ZU
O++V+QRfpYBO2v4uV5iw0Of9j1KTQuhcZSwXf866bJZLGxaN/VDTut8PSAchp/FiCOmJSMPtyoSB
rPs7yGyBicPX3Dfq3Ft1Bm0FWHDEDF/Tb4H4GuF3y0NM1pTkY0jtBuX5fXtwj26LT/pFZyFZjmfq
/wDm3xyduYaOk7GxGE6EGQ3dIQNNfIjG3JVpytmhNEe0kXD5vBAz/ke3OK3bS6kwZ4BoX3f4R/jA
9AYWY/ntJFqYbKLFUyjTN/uaHZEqluNkdCTUZz21ec61InBX1ye2CRymNrnP5MsaXKG51CjndI+M
sshmDVdt7ReWtqv4QNa+hPrGRm7JuQzxkasrM9afA0w/9NM9o3pdp46W/rPahvUHrPtsVY9Kk2Z7
6A48E2uXxR0jytiUjJ37Pl2NN1N+5NoPR1F0mMV0pV79uGsOFSTQmgAEcrr3c8M299x8CgjcLUWF
RJrb5FvrWBSOiVvGU1eHaht5yl3450mXKxDD89ByFSmZulIqeb9r/+yyBeeonKqSzUJZbhYGPL2c
W2Z4zemMjZ8tXqE6TfiFa+seBz+z0VwMwmCrwA6RHB+GwwGENIcXn1nXi3GnnNMnbqcW4YWHWhUT
um/wGOx3hhOvr1MbmygNu9UKRsSkdFc+185DTcfu8lI7kwsFRyyhc5J2uNl+YRgOHNf3amu6YWr/
zSurz51kbQY1/NKCEsWYNqsB3FU0JNIxXrH4fA9zNlx4YcNuEwNPwXunOHg6CwTvlNpIx4RfAdcE
rkz+4xwMNiVw6tH9YiDujzQt6igRn8G9o8QHm/KhtBjXsPfII18xZ6mTts9KlR2nGe++p5keDcpn
AP76zN5aBxSNembQ7dw1Lj6Abbr7I8/QxhbjhSN7WXMjEGOlX6CvpulFmFuUqV480kippBeL/lgU
rLvX1S8KvivjNIID4FcF/Eqxb2Y6vFfdY44Hoh6AxVU6gQkgyiPTiN3sKq7SRwRcqaiGkSJdwJ1O
Z8vnOOrQ6JDZ5iMoGIurBB5y7e/MXV2kNjnGNSPDY3uX2u2n6X28R9IPoaNtkvgFkkV2KjbBaG/D
XRN3lhJWEjjtlxWL5eZMcB/RpLHOYJ61eLMe0nlSXoNUKpNTTRte1Cyrt3Tg2Ug6VgWlWzyk6mIn
uNj+y+vMwzYwVtcUMLDuooG8Fnyt9fjIrnhcR07+aCxmWkCqI9Xh6YVI1Jmb2ULx457riItAW0cm
erxH9z1KbpfnaFdckYGrE3VcPnh0fWiKqmboyg6F98wNStpbDUqeyEIG2r/A54xW+uiIEU4NQy0L
oVT9ziCRJWNrh6g8N2IKRbE+hnHo/FlO4FOP6bgQ6TD3o5GUZtHRXVbG6dRebywBjHKABzxjGRis
GUojgZvd6r/cUcZQcxiQYRiy2PDmtqI//mmdZ7X5kToHWbZ6RaLOQDJPeZUq6dM1x+YzmK2QHgXU
tQMG8cLfVjIzuV+GWp/qn3EXsNdTBDIS31FfsFmizI2OZOoAI7t0MbCfJAVSvXRaZsqDvmdo5zPv
9X7OKYhehRU5M1Of+Z4YxPaMZnUKcN8I54YJtAa0mlSBG5W3+x6v3Hh1DRMCfourYgGkLJuX8yJW
7GGKduGdVuRLsZGHOOHO1dSoERyCrtafzu/9kUNJbefpeXv6ekWEQDDbZjUfnPcwh+0XEX/hXt/A
qlgF0rdQb7iGs4VTznrMSd8MNp2Hh7M7O0M7oQ4OORyfmgdDnscyspHRnMttxP3ZPvj4kIWtxgE7
6HbdC9GOYobg4hjbpHzQ9v7uGJUQKQEWiQaJO9Ic1MX2ZwfvL25gWszm2Vvt55ji/45kK987PRax
cwpLjd7nYNJ2bMWxxCSmUQXEImd0wvRRYUN77JiTe3itLpor57fHhbMzsR0JchBzqt2FYXCJulOY
Z1eLI6rJHBS+AMZv0IOPDVp5KMU3dbyHhaL4+DfLoVzExSWTr1oQboM8fSx7C7w8treG6eQdJoRK
3ZGjZeQLRSzbT88w50fNQuQGjVILVLv2KuHsi3qdqC/MSsjcLOgwt2wdBWQmvcXxJwDM1EaHHbV/
01NJUn9/rxj/B/KfLhVkKvGAmrPu4sGx+pq6sjKGGf2E2q30qF85b9t/YHLLTKUgLI40e4FeSFZ3
LOGyekOP7AtngBxjf9Z1fFMg6li1/42nbxViw2qSyg0ELxE2Rh0PLzWymNi4OOdp+tpPf8ruC2Ce
Vl3cFQnMY9TcT86+n4/pKkg0WaL8+P/lEhVBqV6LQIQIUGmIUyJzzsvewkkPA9OgjR9czcSmePh/
ygUZREBbF3BResBI4AgxaCC+5zTqYCMlLtTC1O4WrQLsm3M96aaohKk5mdN4svD5KTzevtcpAgQ1
9eT4AcmyM9bzOFH71O2RuBhAitS6D/2kzNj76xyySaCd1kTr4qmRp9jm5LMwPJTU2oib9MYRg2j/
BygH7RSJx9Xp4iXV7E6GTwYG3O98osblrboD+EUpMB6tB9ePAPSNoviwtT631a5Idz4wterLf4bA
4esw017QyAt1Hy8X8h2JAxhi6R1o71I+anJYrfUhDSYY5p4gWenuQSuevBAeF5abfXp/sfbA82vb
k1TYINgMGyUNk05PddZiTtYnu7v9c088vJu1dlwClCbGEv34mSztO0DQBdAD4wDLS2MaQZ6taWoJ
Kg18NrIXOagb11uM7rxlVmLudSbKZLpC8mhudW+kfHdnwfFuZt51CpX0z98NKakPKU3gVIc/uIh0
hlcJYeriGFT5Z3DT8aGk48OQr6m+ZrUXu9/e24ae0dOPvRISID/9OByfqifwWElUiFxjnx73M1vB
xRDeHLs4r0NxnRSkS0QWU/EZx56hq5vtkmgdVS8IS2m0sfhoquIOzikWYF1EhnEzkdYNC11eSloT
mux0UX3mCkySzAHU3olR53kRBxhCWClmf9AKoIUV+oHR82ITkpBQu9w+zTIuKYNxNHwXqyKq1cta
jqnQwUIcaVimnPkwL7SWqXW6x5LggtvvrdFWCr/61t6yHORl5GyYW8iHMf1PRKc3XxOaCzQ127SF
KL51V/PCPUQGMNl6an5XKGdTJ/2wLqgieLJRmUc6vBmyshukxxCmZ0lZuaX8umC7AP9XTXQc8Xq2
ih+vSRiBfP3Exj/YpEBAl9tAAjJTegiZC2AF5e1t0sGiiBpFGQPwRrLuo5U5gdIajsMHROh08W5Q
D2fmMNTQvjClZw5z5EYhcr7lIeulcGyYBJu15U4O3XyBNBh+Gj8zRzNTMDsRf6KSUO5W4x3tJ3lv
XpWonjAZWojAwHCFgpQuZSbw4fyZGmQ8danBSWimybm2HJD5+CSqzc8dT413ddqqExDJhdQjhy3O
fYNzbc5ymi5cqjorUCn7G40pLppN1N/fpz3BAWIIrws5dtz0dQ/1PuIqUoVms6IB/A4/rq0WR3sk
ysa9CthcILjQiWDK5fdHy4VB4vtsq+LV0wP69CDTFV5jQuWj+3KHrcI1vVy+4lmOsrLA7JWVeAZ7
06KC+wmAVwKml8i1shrP3MoyLjneLPH0akITxYgbYcI+1QdqJuQ77LoCMLsIgMt+5oP9lU5Lc7va
hD7as8fxVCn7id/TzIZQ8L4WPF67oYCGxWvV/uvkkrgKTFAG17jRlXvNmMGXOlZSMHfuW91+78cR
PkNbBXNQ0RF0MRMPLPh9UtSkRpyi+80rYuUW2RB2V87fFoRF3bKx1ZuqPhkIzzi6x8WcOFRfSKYq
qdSwVV26cnTyVJPmhPI8qAk4R8+b2jpH4xF/DTA7Mk6UgyP+9dXU/6VEQ4QORNL+/XUW4+tIcJGY
I9DFbluzgqRuMnEFxZCyr+GJSGyiI1izewzk6O3w7TFWoO1ueH++9MISvJmoJ5uEZ3v8CUj3Opqi
MusLT8TgO3GFGS55Ed/Zgqh443war22kMswaG+0DEUGJ49Q+ktmwc47jr+Ll9+JHpfTt5qmcZVwh
+GZNZhVSyC2hkcJ9P2yrJDWb/iYlxnCIyHz4Pwj6XEKfRSqLn42nDIVD8zbHmlNmExZ4V8zxjStX
ppmXAtfO2dv0FJ+3GA8uVziQSrnj3uuje0W+uuW4QscCFAQV1zKwn+IkWCglWoZMRE9vZF+AHsXd
D5OvYJwD2vDPCHyXUhoAEGo//g4XOLO3pfwqZg55Q/q8ujtx9tPs9WfffFxgdPlS6Xi2nnrATtr6
RROHF6+L+z+B7PmJhL7ZyCU3OCTYHPWC0axgJnZpEm3wfvY1Zqi0YEfWbusYEaCpF0mfNj/NcYB+
pzDatzhhXSfhowNEvdSWJc7q0HRE3jWjgcxHo+6ot4cqaqq2AvtED3749pABZcFSuOM/+zzUaI7Z
dAGCgjRObi6RbAjwhTBg67NdUvS7bxbWkXPGvIb+9+M+RsclVDr79Hf1Uj2+K0DBMp/EEsl6E9UP
lTVuylLHHNMQmSPYo3XHU2Wd4CHBUtFtiy4sprbjg/ONZDIlqnpb/zmEwaClwmxTrwZmsdSE18TA
nGSbW4/PZcBNh7dZGL0KzFp+4J4rDlrsK7z0+Shi5wXXQFLR2WYYQEbfnDbAKtsT68tk13j+/4sG
/F8QWMb5dxGmFC7pZtNc0683xL8CYGbIhHwP+0R2t1vkwTEJXSpDWnD+/C/3nxuVT31SdrtPLvTS
z3ekLeq/xjQVM8I+cy4I9Xli8e1gBL3sEXLmsEk3kqmPe+8ejD1a4WSvA9Evf4405h+IbAvjcbwr
SESypMTfZEZPiZu2egvbb5sDaTSY1I12mi4lwGTYHoB56Z5OllLaVCoJ95tWQjTzU8THdma9HtYC
orgfPKyMvvmyEH0HGqzh6ZCDuEVAixhKQZncuYOFFElyRF6ZVh+6qIQ5ULKsDzfP706tVfp8w2mu
WifF09SYK9tcrqIajse/nXLAUsZ2zEzeeB+aqEqQE/cWlMKOXFnfTzJXhyofrKc81FLLTe4u1v/J
jcIw1QTPs8zXjjVIRRYKBK1Gvphh0H+e9QXi+8KR3IYfN6OnpWk/Ial+SQnGENJnkUKWYCP+1urV
8nM7gxiS2wQcL5mqazh6Fgts2oA7U/atQw+gY9wMsLJWYdW9rhpfaNTe+dvL4QJfJbtTdbUo4Djg
xfpdJU+jXY5xTr9VIK9BQ78eMvLqXW/sjk61OPebiv3YC5SoIlN7vO04+00HxBZBzBbPEAKFQf+B
20/s2NhovyamyETe5lwh2Dvypu45Ib3KuK+yOPd36k2zM+XAserdhzgDa3lyQlZldmkWtGNhY+pq
Q7NOS2wTGaYiItycImUFkfy6uw0XquXnfbEze1fKjNvxbnAPVYCKBniqfibFdjC4b3WGbO/8CLf3
I2PgFLqoBjyGToDGTJ9a2LgiNVirHFPU55fWS3tYHMMs+AgB89nZdvPbTidZ/Ouq8bIctg6GQZta
5jjIR4d2MUHoCPged0A2nzbGCypGu6rtwtmi93l+LzK9hyH4aS/m1q6i8A/XgIyxhavopXd3FIJI
VSFJDrbjJSM7r5Vv1wigiFhg4pk3yUyiU4MYoMnXjq+TzV5ORub8yI4v9Q6SUC/jX8azVTu3kuls
aPH3IrYTglPkxA1OdTGS6+wRYufguqWbeBCbXwCVtCFkZ/qDILGGosPjeqKJZajZvNJSFwtf/lcQ
m8rT7kCzke1ikRT0sejFIfQiMzHUk46GkIKaZAdUsEXOtRz0PrPwnUlatbXi12VUx/lHkqQ1mUx+
m+IzTRiyn/TloSAEXI0HTqBm3ZnApNswYx/bnBP1Wy+2hB7w9ropuKaNPm8lFjX+rt0k8n86YVFx
Lk00hMCnQqOS8eBERVM3VqnUVSBw+JEax5hxrW2qF5jxAHOPy4KFcAF077BPZ2yO4QzBWkTc7u/m
ktygOunKxDBMpyzvif9FH8djKMmDSDwW+MrVYJIuG12ruPQIhHN+2GSL0x1NBlq2nGV+FygLzGxc
7vmeNBTLISeiumPvdxHcOFmqxeS4fWpvyg6cEpKLdwhMgfkCstsgmTMRWjuq8LIjvt2VdkuHBa64
O3oU9iokWIsvibCC4CBOrQ1k8z7Wd9SO0Sl1d3rxaxOjMf6Bj5SK9+Fs9u1n4utlOtxdclT5lF5S
aDPilrrM0XtoFbH1+IhbD6PCYyXK+Kk6I6X69AbhTTks9CXNeKNh8YpbWa9dQtzq2qidS+W30n22
v9lMWrwDW5twvWuDoO+I0txL4wh5hhrfLh+iI3qeexb7bowWuopfCyXDUUdfJD9NIhjDDOA5yVzp
syOq5w/uf+DTQRLJtzsiBDNh4ZPIy/kBLQ8oTrxZGUnDnYTkGj/gaRVqTgyZFr6b1LGLAWMqWLiw
OXAqVnMAXW5cR/Ef4DWcJ8SNUbbTM0kRHK5Ec63gQs1d8Apy8tx7bIEGBj6HtTVY3SQQksbflgpa
e6pREXoiBxuHHmizTdfs5QzMBszXK4JGNXA1kY9Re/GOP0YjsHkkeEvEVlZwU43apBWxk0gGfWTo
wIcfCwa5W+PUthHJ8gNtsrR9votgDhFAkDR12jDiaQuD/O+QITRdlNvuYhDjTkM+qYIZhIpvv58u
YF7grtkIoGoXCrnT7cDKiR9inFjDmwQt6Ex1xPomKTVXf+PHNIhO93KtEjb+ZNGBqyO8S57EHhE2
hIysYyykb1+fFQbYPVOTOuUM/8KGkSf7vm9pmil81ZN23Clt0eOIJ64ssOW4yQbaMyW1jX/UaboX
FX2wkyKNq5Ez4wIrG7iL1tkC96yIpWVUNJDwk4msZT0k+KKcFHQUsnax+W2fI9A47zdNU2r7Q690
6gNsaJIzF5IDSv/AP/3Xysl0G3GYjtfnR/F0xejVOHY96JB8DkJ+vyExvoIXjmjmVbnWpGdCg0IX
G3SZ71+GCS9A8hzjV2fGY0gVV6nHjiJrk33Mq9z/C5gyS8VduGo3dF++VYgVdN37zYfO3ev3Qg2H
WreCdfVWcVjHYt0QXToMWq5YAo70sPhtMmnH3dlnaUilZw1NpWevIIdodoJvEa+Xo5gDrcb6A11g
8FKbdl7DNZF06of44S2QeBlTd8rkecw0QS3BvaFemn57zqigI/8rQ8QLh34wr5Cf1nQaJZVqDa9R
aWyQeZwCDAp/bnNIZubElPhQYAf5+SDnUXRx6tv15Oe+7r3Cmy8w8u/8nyzBNiMSEQQl97dH1QR1
9vAGA80bj4uZBlXPdtProx/sjRzvv8lIzxb/VIWfE561HIvTn6znpqRk0wqVVDrRuY8+OA1d1Eyt
kx/Ah26G+5iOYkXTcIA6JZTu+6tE1d81gIvRFYl+jPUUuun2hGHhNauwJg89yRWhHzac4w0vvdnJ
Ha7VW7amm9Fi2hBMPFRqcHkAmDhFgkWnw3YXr7fbQZ/Jt/DvZNWD2EyZECz7VojNeW7gAnR2KsGy
7leX5mUDZbnhKUmHfXjmAtIcB47cL1twDheYG+rNj202zkHj1dwD4Pos3vZ89eJzjsEgWP8QOXIX
krOADY9TXHDIAGUUvr3BctLe7TR7gkHaWzQ8RfPzUP9lTkhdaeN0+HvRAN/Bt4Vp/JndEDDwPffC
C+4Wn4Dx5fCn2of93HwzU++D7SrePamaiMer1T9Xarm+LbdthySPElEvDZcAL5LNMOqPSH0rt65N
d7HoJ7CYrbr88X+4QOkAEcDrsdxE1rf88GN4yYPfjhbglM4Pyo3/CHhJuhcWiDEl9OC+eovJS1kK
RUwZIHRgcOhrmAxHJ6AOnfXktJGih791kRaHjVH6SZrRb16SFwtRnDkne1e544IQn0Z0/1VMU50O
eJ2x5CWkJxOT5kY=
`protect end_protected
