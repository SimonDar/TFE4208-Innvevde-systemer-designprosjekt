-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Iqz68X8fsdk4RarZgtBNvpW7kdUqZLHUuW8ta7ByOtvJLpE6+0JGdJiLAS28tOAlU9tahYYwFZtf
gt0msUNk6uufllUq2v3qZAQRpZQt1ZGW1tynhRGsZyNGCXEDc/FieUKNg3S2EcEQX4FDNluIwY+D
N/SZe9vEBNxL/1+kVzzz5bN+kzcdpgQz6L5N5s4MVPyEeEHm7jECC6Efiix2+73yMKkAZeDWZjsO
koOXMwe+tBW5rVjMVK1nimuZIfXrkvZhN86j1zH2CAMZIVULahflXO8v4aP+kQrOggra8ZNDwk0O
teRwEzKN/d8ugiND8JrUV+cQVhQTIBdqE0Lp9A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
+JTsiPe7sqEvlBFxx865yBucbwFs8lcCfuX72Qm6QzbtrBRDglFI9D4rHgMNp/8CRo0veP+COcy5
wW/3hwWgFnhERA/YCSv97Q0kPn42oqAnFW/oe4V2wFkTazoBdBifxmHExYt3htZPmjt40Ur4nKrF
EqWiEZyq1BoMmxLD71hm7xBrFRtjVxc+sn7ZWzz6r/5CDlpKHlvQfb9ncsaPnuyNitS3NxKbcu6s
wGrENUUY23br2qgPO0KjQvDH8vZhGKptK4nRCka2WkW/HPMUnljqS6QzyUP8RQRMytvp+rr4NO/T
jwaE1amsgbT3JX9Ji8kTTb/IRAqt8gqAKZf95Mnjd1iBsbkAfxvTIbKsEQ2EW40UGaoRqnsF26Dc
1rNeIJffrNeXyyda5ovrFL5Hyq20i7cscVU8D6PfpmOml1dh512f+nWqpMjzLf16iqSN/f34IYd1
PQIKptXPBjQVejTNHNnJhQg2mVmugcHioBp2D+RbtVHp+5w8d+f5Xw/ET9lIM5IhWFL/ZSdS2Tc1
VJCXdyAbV6xrWkIJMcsVm6z35iLhC+5lXM//M7AQGPIsmE30LQbw4DeQB6xtVzdi9fohj41ZeLik
VQ9WeLMtERaJC7VeG+4MKbkqLVeiLZKDBXTzlsBClpbT8uCrV+Y4ewDYybIW1PihI9v7xmI46N3H
ezBiuIAQgTwkOly6WScx2sQTCphQGirPBCs8a3idP2lst66HOtKstt4ohIFJ6SKIz4VBaaPR5P0H
BFNnHnEPj/nxsqpzFV94w1Bp6ej9TKG3XDBm2UV0hDmTclsyp1GrCEHDX/xwVFcBQaT7vBPqbQmr
v2UgMb1KG4DKhXNE4x+/g/DlNZkISka8VBZRzKmOMScFXjlcBtmihdgarH5vxnpbZ+KG9jfj/Tkp
BtjImyX6RQr/RdgdlTzA2DmMfleP6mAk/jl9LvYLALu5f/X9IaLBxha8HQaDZmEu5CkxffNw1Wik
Z+/tJH3M2KzPv2TsiabYeSmXDoEdtqI3kiGMogx1fpmYN7roaSFdi//qPbH1t4fas9YhKcqVkfSY
CHadWbhWQc0K/ju/8VzZCTXC6xPshfjvjhj7ZcQwkvwDOtPETEUQbKfXhrpUGXwOclUC0Gq2qEJR
5Pdt9a7kLdOgXqUnnrEKx8NMB0VOommQwk0bsc9VyPd+7nHnsl4IHQ56FR484ChQmyJQTSZ8JArA
oxo1SuV2MLiaV1dfut2pOXQO8y0J69aWW1prmByTtcfOnvuq2chp15v9WO8meHA3jO8/eMhCRRkc
Ei4lyU4kf1e6J1LoU4DWYvHh2VozrbOTcTLQHZPm01LrDNL1RDhr6u3YBqeOPkjyOVdJrnzIZ1NX
o03xvCVmfSnboY2EZZjTGO8+lu76ly7Z/cPBF18KdUX7lLW0pO/Y480miY+APB/9j+l5dTBbGUvJ
g8IhEknki6Lv4dy+JaD0/Ndkd5FTc6KXDuMKl8gVMxlWJrV//f2DMNMuzzcCpEqUjboVq4SQTGVg
v2Nnj0mKiWQ4FMg+ZcEpXZpIgj1Sxe+BWUFewXo3eKt9lQ8aWTFfwAnkzslXni8nwmxnXd4Ccni6
4q9+/PQAa4pw7EmUxGPMr1l7zOE3aAN7IjxJt9ZpZi4lA3dKeTQfcuyNwzNfjwNb+nrB3WPtUXay
6hOUmXLO4st4Y3fbvGf5BVD/QgNhgRqK0NUQvozqwV6If5mqGZQVayWkqFPCPT1/+gB2ZrkOxYA2
QImxLxy1NKE/2xTMMHNolMqjp8v74wTdT+4tMbgyRic4QFEPfdMu0Dgc4jdgp2nhv4KO1Fw3vK/t
PSLatr92BTji1hyFKrEObundjPQYkPU6xv8/5ssrkRr/uSfYAzKimNvtZPeC4ZwGt7kXUYODGBw9
aF26H1IH0qnpoi0WhIZ+uGlkkf1bO/yzRszrfsVxhbmBflFtsX66TiLDy/zvtgsri5UqJ/iRaZyd
EMYjEEiQhWfrt9KT4jRBuOecJO8nMI9iaBIziKv3/ugypN9AuF0JycOpB16LS9i6jr3mDHfiaduP
VX64ZnKVnNZWMqpLz3ZWymnmou6Hie4i/qOx4VdeFUfkxIY1VQc+oVEH21WXN+sRN2qTY+R23CTZ
saK6IVrcJZ3QKpq7teomRGabsLX2ubl0/04YjOJquxcaBFvYob2wKjojdU9oNmpw6QZB09yDekmj
N47tHyfqMCb+y+bmUO4VaEEIT+Mt/lj1bP75m1vWVpo/JBdurFKJbzRQRVnuQUQrrmxNmtbjKylu
q9BNnbjqeGwshp9Z2pvf+AbkwuLVLPSrtVpHIRq8q85aVUzKwlNRfh/crRJXKRjeFaWwwtyQVNfm
QQt/awNLJVAiBFD8nmx9oCb/8aM3Bv43WzgqVNu8rqJMM69fYi8v+qza9WQHSDxrcYfPdMEb9/P3
Z5qXzPXElSwSB6f76K+ekzlU8Z2r1m7ob3lBgMPeuxnLtJvu3/6t3qce62qMUeQ7cSHdj9qnEO6H
jJbPz8BXUCWcgCaGKiNpSqAW+DefTJ/Xmo7Xl/tKIRLZDS4x/bcZ4zFFMtJ7gupAqc0NSmbw5dsR
x/74hl0qo3x6KwHD3skC7QWRwGS7sgwKtYlqS1hk+Rlc3qYXkYszOQlTPLma4GEFJKlirMZOkT0W
J25GzHLX+ku0zDJqhh0/MYYJiT0KEG8hMYRlAz1Qtri02mpMLujxItirwq9+i0Y1xmyfABFjBkcP
3C9VZJhMASd7+mytc1NfZe82D+0LwoKeM70tSsCrCDrWsjn4vAs9TsfzhAeAdN6khT6xOkoYPWW0
8sETdOEb+07W9XYh7pmXBW6jyOONzeL75wXDJy3ggf1jUcAz8+DXRXpU2XMiMfMny6ihnGbAn7X0
8IgNLPbpNuIZglSqkhLFozXqgYY5lQcRenTMOglaKdy1Tg7ngQ5O7KV0trAstyAfTjmrRdKr7CZY
hpiLNkA6JhkX4trMph7TheTInFpZENZt851NvHg8PYx0+bkURHKPyQBOjprKzwKPIvguEyqFtNIG
6+cX9QmUYY3964qyM/WwrEjztdXKEDcW8ZLagLO44qAG1+0+oPyEuYo6PcRehgfgvItfyJYzNuuc
cP/g1yp5ibSFyCz+ZAsWxxtGhUiAFDujSVJs6PByIQpaUfEM4mGPK0WCMugDjUljrE7AuJwHQARa
npCwbVgLiN/gfU9XmbUKJwfgoboQ0jLRs6iGwPoDIjTlLzXEwZ6UpqhERUhxx3q2GFmsNMVKpVkc
Qqx/pvqY6HYA25y/5XPN7GPEHFu5ASOOTiPfCVSPt6WAeHVNOl/TRT8BZADU640fHi45IjkB0Y+J
NqjI0wv+dBlikC6W3Oj0Ie0hC04CC1/UpOvoNwkes63PMrZ1xe6ou7CkPkub5J4eMnfiogDLk1tJ
dXY0NWyrKEhKlvf/NiEh4516JWd+Ncwg42c60+uBPPXfYecybYSaoeYjNyZORMBj06GOE+KtgNuo
EPs7XoAiQsXNWq9iG/VZsSH5sKF/MdNKiX69dU46P7cwvT4IgyJmpmt450jClWD962Z102tw9zp/
n5uqc7Z9Ngw9JZRV6MGEkfu1DtBXYPEyEUVICFuxGaSu1woz099F3TsBN0HnWN0o9c8De2O/1OL5
VkZmloJjs/TGaf9YiV0FyZp6AuU+fCip4rZrIOc+i1sNf4tzHX5EK++/9HpA35DjgLFmuZgNa16k
4Vjs2L7bVlzyxfavUlICacXHSUVbtdc2i5fMSfGtLGkc8UaKpXY57dfhDg/ExTD+gAZW3l0AVlBN
B+cmRCv63Enk8kmB/QKnTHHWEWEbOYLU4dA0OJUgrhIKGXm7zxRTb4Bn1NprOw3sSIjMddGE2MaK
tMYNiUxUHZ/ALkra4c22yC3f20QTzZErI+ShS9aDW35dBuoNG5hwrXAW3vpC2fz52XzkiUpIGz6i
+47vWfZewrkxl0wk0m7G2Kp8wzcfsLr/N5IdIOu5wXexlHbDnJWlYtGE9eTkcqCUQhzggYlT7vfI
QSzQmXwV8oJKGFakIRDgskfeQmaFD/iCznNwMK4T/8Hbi6ozI8MER3Pd6WVkBK/fE2I0GHFLUfui
VSK0jAkn3zzDBbUNk9XOYxZOPHl8XUDXZJkWKd5s2I6ygaQPlJ7nxKNPqs7B7RnjQNAspXNgtUVl
Ymd1tNlGbfEodHl7A7fQDaXsQo9lE8CGQIicc2/Y7WApR+LckZqfUnoZKVk/gxb4nHSk505DGqxj
SnxEcN6WSSg8U0wi0MrN07d/OcGGZLU2rAdY0s66U6WIMEG8IaMGKFSbVJDcOhId57ol7+J3g1kr
GwAGg83Xqrd98ikSXhQRloHl+f7BEsSybWokC7oD27dmHpWn5w5WI7q6mfY8W6CZwwOP7fo5mHgi
FgJA+ZRP5fML3+durZCZLhGT4IJYNL7ZpLVcxWZwth3bC8g6LHN024WGCt37Op6Nh46oHCfGJI8D
+0GClaY3tqJ/bWtmrWrbCLOPVvvyiFsqmGFWxFzfbpuuT5XRXXMRnd6kPwoCnRLqjusuJyc0Rj+y
1/z//J9SzNyOTTqKMohuKxVEpNTIohtupK6L5m2SBRAJl5Hhhzdz6ofdivDqQ8usj9ETR1rjcvNe
jbXdS4cUlnHKmAQMB/XQhAGQOaq2BFIdm+/rC9P3G9o+uTWf/DDQ938q+HeCAmRjiUgyAtvy/h/I
k0ZfngO+Y7V2Ids8dtAX1IiUgJX2fMELovz5R7N/uFv8j3pkKpLun1wn6YPNOdRnTHXrg6VnAtar
L1bBmg4X6alBzUM2m6w8R0FurrGdAFo9oNSAcyoyNQ66XoPmn8slYCZDTNo4bjG+rl+AAfDtUK9r
7wF+AfjZGx49eMRw3yaPhbhYrxDANlkpdEEKTXtlBJ0NaQcTvFlpnXUIrmw9DmEG5PoNbdM8aGlx
Hun2V9L1eY2vWDzYdd2ZeA45nzHHBpXqbYwd1aB1T7txqbBlMeXkIxM1L4qss+aZgK242AvhW8R+
eZUhoHf2HAuoWc7pbLp7hsblpITPVObRaynWRMS7ac7/wesxRdDiC57Uy8M9eW7Un0Fd7aqJrn8b
JNAGXEivEEIDtYtkCj8Sa7fJG16WEQoGFCs5TcVf+5+kwVP1aXeiEE+6pjtaOWP69aDORueEs1zH
425k8//sx/GbCETXy8JS3SMZHS2/n8ojwvX0OS0Iluw6Vap5zMmsRhaJi5M3SoTXtVPzBGJEEEG1
ID5h0TMA6K84tmymVRgOR/R3NIJ6T3rH88hODzYNkI/PThnMSXq9yZkC0BlCtr4b6fVRuzfiO+tg
1bu7Fpx7xEdcNVUOc8dDE1X5fHZpzlZhND/I7XBqYa9jXRbbLz1QAdkO3PZQiEuAq5BKeZyHI/nu
unEmnFXM0RL1a2BsIDVW/nh34oPdzZ/LG2KrH2ZD92Ud/xi4f+Xye20laDl0TUDq7DH9lY5bQeEm
r6tf0l1tlB6PxRJNX+LVbrNwD+S1ZEMmPgR5+PNSSTo89iDXt+B7PTAZDhZGu/dYYns02lshICtd
nuxDwZjVwTzmfmrS4UcfwnbvCfLSUeW6Y6BhWe43GJwQZaPoNCtWYptodVs0nzBVhmGC9FTpbmmU
osOgxCkY4rPhOZVBXvJYX2tdoTzSueU1iKjqp54WNoBtE1namZC6DxjYOs41Z1NCb5tVd+sinvsJ
SXsDtZXt9aNa0j4DS9dnGtdqwlIMWz0qyF8uYir+MQW6SlynKa+fVbxp7EqnV8BSfpaVFi3HPQUE
9CH9NKiPX8/yrrB8repc702A1AiWV+HxAceSaAtPJU1+69lhj9lUeaYjFAzQoKK/QiiD/jhFHzxl
d5Lo9v/woHQxP84LKFQnaalwWYGwFr3rRVj4BzKNi92BFRamCBucpOGHJQzhbU5d1iCHGuZwqu+d
2AGnCD0omRyQya3qmue5y1XoaN9a26BntMOh5DDtiMSiitD7q/TSIfyRtGjaXDGyg+fs7/HMdy6x
Ti9Iq0eB80qWZ/TYA58OYgvpZPgb4EgOCGa0d+AlTlcrJDAyiX/EX0iKk/tiWPk2aozV+UDcMeL0
tI8WIwloBJLYYOOQKfhaOYixcKZxULs2GFmTa5XN+zpa1txHCUYLZ1efX7hdmVOp1GICAEBoQ+lR
rpovndz1cZqZsRiS/JlGd94wj0WAyaIJjwkmA34FnJlsWXDNZK3EC4H0Vqrpj+yBChce5zv1uDp+
GJFQRJDWF2rjn8UFYstXPR0F9iy4uZYROUTsB5xckp2RPVbo8pLHLb9rgPXWFCUZGaT0kATPuBwh
v3pZ+lOG0w15aWORXfyaRAivXIKDEE0AXljuQYv3aRwwxXwQhMTUKImYhUjpIxl9H6bDTvxREq1U
XndIMuOA5CT13CnHE1v4Hsdbu3XrY2WNPDZ/9Of4cLHij7o618pcvekXr6uFAYvmZTbAuADRFfyg
kLjBVgde9YsIgvmh1wKJtJj4klFfWD6DbwRvcIp7ssQeZ4Z1HSYHE41h3YSrDQrROv22v5GxqLOE
cvoMfmPu6kKVu0AUXcE9YN9eoq7ayH8DBLejbnTnfo+biBdD/yCPM/AFD8TvAwN5TFwIN6iWUMkN
RJ+L/1xYHK9FTAtRFzjREKtEXKWkh53f/iZttzOHTSnIvRB+Ox9gbW+aCUkchXvFaRf9D5HD6hox
/PVSnCLHGqtGFdidY2yA3/QrK/r8JXexoCTmL/xDR3zr3cxu4qzKptPDdaxdv6ef/ba66tIb2S8o
22gxktlP5bEZqCYnZjgRrEqho3v6WfrFcQpAELYBXHpHzWsiN2fykJNQDBo8Zjx9MICJ3xGQaF8S
+AVfZ0LcVb6EUfwC6KV6lNW1IWc3xRV7bHNxH0Q5tCkJQp53fEhJM15KY4b+Tdiq/0Crs77cxcw3
GnbOA3Ct4ZmTU58JpPokze5NTj8qpB50SMLWvWYVn+yaDqsojL6dU563TfZGkWo6TyeckgazNP6f
uGNtX2l8LRGtxl8iNah6LmfsKELA7Q/QNRi6yRY6tG8jXlovVCyiqo+HTeBXW3mcI39J9h1MtwND
ZOssXTti8sDPqIHFXSXtqJNKKlV/sOssFJpYn+VQqjNsMm5rUJjM4/csMIM3x1kpAhsPvEfHjIb4
160e4wlcTWf0HMjMMrSV+fRBlIROkKZwiQ0sw/GcTUyKU2USdYE64ydOhad8tE/zZ7cldnnT8jn0
729TK8tug6gnY/yhIxM56jmwkvhV53VS07/Shrj1NJjRo7ADeC7Lsu+9RhOsPpyJLDjgXK8Fqga8
6uL/HAU/K54c4NZcpyQ9UEy6IR7b+QpVudX2Jpx/IlAY4WhuEYxdhAaFmKLIalSHxq95ETNcOxU6
DxMUd7AJ+CPqk95wXdJ0m4ZuvFN1/KH/THiwcbhaeWmbmUTyIqdEx5Jickzzk0nqjuX4e8fb+Wok
hq1IeOhyHT18gx7U9MmjA4xIWC3BeYtiJFICGH4JfWb/S6ruEkoS5dZrmn6+eb0leTZYMBgDtB6G
COoyo+YShyE/nj25fvVPkRb1lxxp8VXQjGXzrHeyUpL2q+3E1RiN488W20qG2+N0YlIqgzD55V0K
CCWJuOsb0/QcvUPMsD4tU/lgDPUWke61UbsSdtV8ZIti/aWU+DDht9I6btBXkilFuLDB/JxrdERf
BV1FeuJCkx6yN8COX73GFchpxHJYW2qQzSu8pNsSvKtP/2otxpECS4S3NUJOPCWQ55bvIb6cxe99
Dkz7Oe5fTPcvMLkyp7RJDYQ7YEjWdAKsfy4ackyqVhncAlvs/h1h24e1JsVl3//OIZnXMHPw4Ojt
Leu+NUQ3O03DKw9Qv0zQLb5D+jbAsQiMoHx86QJzw6/p3z/SeCIYGOz69q2X5p/BH9kfCrv/5CAQ
pbhJFkyLOkF9PJMyJTY/GN0i9EW2HFXRCfl6QmC6eNjalRhKI9OcvqwTm7T3hMzldMV4RYeozCf4
GGT9PUcOCNm8n2bvRMQbVAZjjrjdKryKsBF/nV9dtPYaOSV4MTYqG/SoVEVl9TkOU4QauQzVKxRf
tL6iQ73FGWvO6EFA/Ag7AJRNK9Nb/y/dtIQbMeQ2IvE886uhNaAaj/3sTtyt8IfaiagGd7Pi4r35
wtlTkspcWAfDjMHgMNXWS4FAYkT+AeQO3hrfv5kv10vTVVDNYLUxr3tjlkOza1CbVnZ9Aj5Manjv
g3+ufqY5EOH5r3eZyEq78nMS00a4s1oohDSp0Blh4QzT51XBFqyJJ1+vS4RziF7mrZtZ7DEUTb9w
ltCbbnLqfz0gCXpTqGp77FnVZEM39/SPWNwCCuJa99hUssq1pW8zbgRbm2hq/waPm393OxCPl+EB
VnbK69D3E8nofB28oueKiXuKTNNqvk9USuJGWyRGfewCfJXqkJC7x4+18QPA3hDPsZq1lFpArwUq
2FuWkK3Ebf606QzL8xVfJFpduJGFZ2UihaVN+mbobP/3w+N7qkXETVvbwetSjiDznTjqJH13PHQL
5JaL7af9IqZPRpF6/pkeoPboEyHJs5lIrQ8GUyVAHy9CCQwtTT5YiCbJPqwt1juAPKMdREQt+bZq
qT29PRJH3MIi4AzE7EqMCTvsZBAm5nyr/CcAc2b/Z/0v/62HaWFKjiD7wSurw/b17+QZ70Ihr8fV
i9oaLkjLBGPxXwNMG3xV+bGv/baOTfUYC1Z+izaIF6tIk/VGXmImNRJ1KGS8CrLDGC7TAJ5J1ol4
pHsdgWeN9Etx/8+amACXjVAeJ8XNu1aKYbako0S4wI3awAaydvBaFSyIl/JyKtwxyJbd6MzSEQZu
5fNEEa+gEIKabPodlVpTFCpNv1UVGIWFk8DVOU8O5HA6zU27PPxMPNFlA3G80tYJWEkXxtq5PS4+
s+yS3K6f6VQCjX3Yi3+3cpeCmhLAhzj8tZetFpGeutcHPz+5Ty4UdxeRi3N4D8TPQoR11jBKHnda
LUAlr6+s3AzFpUaaGo3r/+xiUGv5XQ9drja4bt5cvvyOYnRlWW2BJdBdl3Ld/zkNxwCUkkjFkAXU
xqG+yq3fdN4+yLjIRm52qQqk5FCr5lA1FzSyictqLIJ1+lON28/P1JU+uS1kfpkzz8S7CWhA7376
Cn0MCFayTxvW08DAh24IfR1pc57M6YimjAUoPOrwt5vRoou/15QchNHW0dhwO1PWnp9uQOG5leHP
xI6eNIUbcygCqiC++Gnphvd0GMmBbCw37lCcEFvnrvnI90o2hjNAkkCesfE4azYcQIhFqvF8gZc2
zzFb542V7kGC/7Y/v+Fgfvtuy4OKGfAA10K2ljdG2KI9if/jVgO128vhCVudLmKgkLeJfeNtOsIx
ik6mzIgRtVCibfwHf0MzRcSDA1YcFoe8+2l43GEnTxOOkleZ/B79YxpozM7mN2riiJTNKyBlVNr/
+e5oPynmQGpuppuGq7KXn7yVjtZ2Th0r2He41oZ3BPWB1ifkc/kTfm9er8E0/XuhVy2gGFrIjCNN
m8flWasgOadiKH5MHfaaMkGWL6jiwRxTdoHukqRPuqOo2V7KbpTkDU/gPr5WzoHcbcYREdAINAqF
UJyiqvapCSp+kBAdpcI1l2VutbIOoggr1sDQ4KjVsxZn2dU9yKRvjMf63OwHp2DGNksUeJIkuPG6
l2ErzfsztbquOu/7vnxomCx5KSTNcK0JiOvprNvoeQZhOCz7/K0bVXHJCQe5yYzImV9PhhRpH/kH
C2oiCA8gC5khRF+IkQgmohr/PkC4TDTnXEdbDCLHm9vQa9YhrPBhNdNTIFY3ZF5VDHjHuZ66Hj5U
S+65xvB3uvv65MsZ3Bj5oK51p8EvW1xor5U/5XbZOFmmMjep6Wy2Za2FZJlCWYp7W/jaA0txAxcI
IDcqiQQ2WiJ6xoON0ytMmY1P2/XudbWU8BoaK17Q99JWXpvZJzt0Xgqcf2if3MkgKqw3uFO8z6Kd
2Vv9bb/zabY2pvGisRR//9wU7oLANHSue9Dncg+XKMhRpgPcykd4H3woS7kA0doqNEooq4QpVouJ
Wu/r9D5xNhO2AyeYNLLNB5zEj0cZEoDwSPPioK8My8IrtG7cd6gUA+yEZMcO1fEEs5+aBfiPcKNe
ITQNXSHcUDpRTktf+ivtlyyWbQiqOqPiCtx0i1g1WRwdm/AWb4qp+1zfRcF+bFwyhB1Q1rx2cMi7
Ugez7jLfuNZz5WbMTT3YuQ1YotWOa+tnkaADn1nSW0/cN6RKZLESt1LOJpXcrm6zt3YFrjiCstom
HPGEj2CSfAIgcAMNDZByvO9yldDs9HCOHj1h9CzOBPyvV1wXRejPFu52n987GC+6D2lDezJ7IxMR
fPXuNZtvjynhw9hNBCT1RPW0D797QTfxrMa4DS44nMAuPlmTuJ+q+1Xqk69lYENh4ylfEUpoINaG
V9laYqpj1sEQDZM7xIDhqYFYjOSdlBQNJFTqqZnPOnrQrvwvylmIb7MIhGj5ECF46gVNRLDabPkb
BtOMxBtOrbwjtx0NXk0k2AR/u8MklRUy4sVc4mzOHG75KPzp+g10/0baiA+ETEqTjzGKAwrFVhTk
o3VmbH542a3Q/niTxxGSmRxB6XUdvvRB94GKIh8IegWpU4hSqN6Yyl16ue08P7Gs8lzwUJoMJcRx
uMSXaeDl+fiTfWZHxyQbjBqwb6fpV9PDIYAyY0THjLDzy0vJ9MATPs7rYAWE29GrktUUoIrFHraJ
zj53HCkkN6HAHcnXgFKvd4DfgiCDSBcznasyhsc0wmbjwRgowX16G4GrcOBIDcwNzphp/GpaTA1R
ZU8hvUHE0m6tz33QFLQ3Ty0X9T+piihswNJM25jY6kJuKPJQ46dTDDGvNLXWo3bJj1pMCFgRjO2p
sire2z82elkW9p5vlsi7uqcyFxTSUBs87fNLjL5hcfj/hkC4PChq/tJCof6xBYPU2sRPFPXpyEb+
hiZL3siCTjCCE8Hlf4uHFbX7fHSdUXiqbHKM14VA51/y0r7IG3Vd8YFiR1NNK57fYQGUxZr3rbpA
aJ7VAmzmhfg4/vw19YOY7aVEkg9elqd4+5WjxDrEbJ89UkNX2/AYfKB4GxMWFyw6vfI2hPJjP/a7
GhvUqg1/dL2Mj9pZKYPGdbIz3rfToSmKBwjI7ID17RCkxwm1fBv8i2eOVulwuvBTc509WSCZN5Uf
gTqMW21Ib2v2CkR3xHaKdW1phlAj7SKaek3roPoHnW4K7ZvsXH4Xkypux+SoUseqRNRSxsQDlMYA
nBr6lxN2YiQng+E591x7iM9aWxcLPTk6Bb7qgAfNgry92Wxus9AUBpz4GE/7vpn1y0LHnJWJYWxa
dcCpB0SBo4MG2jfFC7mCyE7cC0TFL0jaJn7FC4/vjSIWmr36KNtKmIIwUx4DbM4cCkkjo2Bwi5zp
g2jH66ChBx/M+qlXafroM2RGQlDAar8kwEM+IkF8U0GXqvWNa8a60TR4y2rkf3hgt5uQqt1AtXie
Hyu/G/Y5dtdQBNaQS/2emQ2Iwdo00IwmyA6io4TrLaY2jV8X1fHTNdUfm4zeTKW171v/0aWKmf29
3HX193Z1pMZVNhbvESh6yYi+hfy2+2G1l2IOaKZ70NmWwnQhHNVPXSalax1xc+Y4WMFVH/St42x/
PxZ6c19IwlhbBgITFlEqKoYcQcQRoQAXB4RRSr+USfgqxQF6nN0E4DCVFwhKgl7Lk3Xw4+4hILeZ
bOF2UU42bm4prPPldEpicCgAd7ylSsPW1UL8nHlAOpTkPe5cS+6z42DLagh6lTEwlbN6PBx6c8Gc
MsCm2SEhWFOvYbsMyyHAQnRiB7PK2mbnkkDajEKlC3Kjn+XZ1uckugPQOpcIrT5R8ZIyyGQgBf5r
6HPQFrvbXwsmOLAT1QzuO2gsUPD3TN8acOjChrD23n04kY4yK/n6IvIlNKaO3FjK7ayo3ejqngk6
nnRRc3NU2G5SNIO8t9n/htLW+n/Vu+Ws3tEYBvpgAZEyQmjH/K/KPuMioUEf3SQ7nC3SC6Q8TXPw
T4SPZ7mEMAbotxHIkLot+1WBtpfcOZX6UQUYObYw3e3/2TA2DhLsFQ3U9GxB0YbAn34lMH63mDY4
7ibXRuKjMxEd2sFgJ3oaE8jdS5ZIu8NJzjlJwCSuwCVT/QnmYTKB4AgBqbp+a70hi6P/rvO8KpZQ
xDk7ErVGLKra9LgSsWW4fo/mX4EVd3W6uoYV5fOPYxvB69SfIuBNWEO9Eq6+5xPgZItOQnHWyuJS
p5oeiwQiYXjwR9euf+YHQE2EwB6CJuMdH9A0wz8xY0AtEQkrrStKpPKCt0+u8gv5DLLUTPxCuxiN
gkq1oMMOtaziTVY/J2LEtmqcKj5XnHPl5ElKJ9d3AhKzM9L0x+gKF9j1hG/CJEWXsIGClG0z4LDA
WTo2127dkFYEvNiRnDqyltlNShDJ4XjoEqXZtJzrY70yg58f6MUA/DqWHWxLRCUpctGGFYBHVPVL
C5lvBebwJmUwRADdYAIGqrmQCXvYKBck6JyGNp+lRiCw+ofe5GaJixoGvcXPWfFeRTVDKGCjICAq
gzJnNCo5j/vZGOhBk7f/RELyeHubrLiNMWbopN7ktS7DvSvwoi1uX65MiOVEHGaqK4fgMYRddHlr
hcrHVFTjd1LOdF5lS51r6t17KcA43KBFlQe3H1Uifmw1hKhUIjZHc7XD8Z0tfnTOZFsFbYcPsKHb
xhVp19x/S2PgQLP0blZzAWKga+toB+OMGDSrlM4aDNfCxX+LlPbEH7CJuZ9CO901mY0aH8+r4R4d
/hHUKpyclIGnnzblNnkGq+P7dZINP8s0s8hF81w1T9tJusVmny6FN4h1nSuzNn3+VzAIlDpgwiME
ZR9zyI+WPNR0WSNYdlMeKZaC3ivL+Mxu0KcLGUVm1DwfP9A1m3TIMvc2yt3pbI1VZn8GFZLoQjCZ
08TWl5YG7lNrapPppg1LHNUpTkg0N8nugHUru0AmYUPFfdAy+HSEOjqNvQsBcL9Eus3PAKuvSUi/
jugaXy2Gsmi4L1CI056K8hkmJNSPCkkglE6jpHjB3f2XXXldf1aWpTBRYYUBn0eY+KpjirT8DhgP
Piv3duoDsQfOwKbPybVgQu++KFEW9x9W0/5ifYW4mnnkVRhWeyrIfpzWYSsT6FT1kDcyPI216aAj
FhtkeKCMwO+9yLS7rAIvBZD+PrLvrIWOTfR4GcQa/TnkeIbpxkh4e+nmuw7gLmiGPBGYXr6U8AkG
RNwdQZSJdjFYl7xKLNPYzS+vZW29cI7FySf0tGLlmLThYCHTL7x+ef0FqNFsvdr3imJOaO4suAs0
BNFBg6H3av3za1jQBBirhGRH9zQKV3VfJ8OvJHLGjANYcv7tISr1/3FIkFNWCuhaLxKWzEeoSOaY
/B0c4UXmROpD5E2Dgd8u+ixrM0LmWcqpmGXH0BErxz1xLwyS3WQcP17VqTtFxEd2VwaHsUuSoLHd
NMfOLE774QrvVWualRI3ZbdaykS9ODVgVmPI5micRx9CYpEFMkr3qczmUhJe8AuLLPxRD7w9dlRt
ODHOG/wpRhS38PSuRcmgVgnGdbIBEa9sKM+gAguapwmv9OEK8cyCRMlrVCDTkH92qr3FVH4UY2/7
FWjF7OIfw4zhBUkyOij00ThsBXp+gl++uJuXN3Ys632mG9FsO5J9pI26oDUHQP9tcccjmjU/YSls
T17M4UN0vh2BilGDZnJvQ7OPR98MSCfrwvTFMqY0AQMsFiVyaFuO4NJgyq8ulwavzIDyGN3t7QaB
pT+/Oz2GQInvo3PMPyHmX5JCzFLsDm7MDP0ibh1wB8zRGwbF6hsCkRnvCD51Hsu2H+0JvFM6K+vX
pDzAHyS8gY66z1Q3hq6iOwr9FhHvxUlUg+mu05ZKMryz/mZtrZuq+sF9kO7dWu555BxQnVCWvgxV
wQyAGJj22cIntyfGVJhfgsNUc71TOKf9Law9aF7Qs6Ns7Up6xWieOstWzYr+4Kh10jD/60ylCc1L
Ec/gBszILznhmjFbuuXJIOvZItA6UOJBtS35Vf9gwV9vF6eB9vvVGD6xXD02k6Co86WDVCRhkrCd
F22VQ7Tjtq6nAcKhntJIMQ3JYuc/JAHc0iHZPY+YGvdaGdXJ33ChodxK6rnuu1wS2J8IhZFsN51t
tGnL0nY9gvMDqOBVHMUni/uM7SQxep9cxkgcNArPcF+o4te51VwUUUyflwJfuOZ75moXDSMlSELA
Tqg6bK9Mqd9Fwci+ydm66o111e9DNlllIjsyVeSR2WeXK4ysFKVll1c8dU4qJc9oBZGTuGkYfXof
VwHIkw+CUJPsm2oslQYM5TlIkXl7NKbelalDwZ/NO99+eADaE+jTyxGepJbPKhTHNLuKWqzll1Sk
6VIbbOIrELPxTy9iO21f7BnvLmhgYtuLFonuzmx+yx9NPfg8EFHaxfaCEXVy2xyt+ukVERtKK7ng
dwVEzGZH4OeuMFLtxBnArWHaQTumAuRnNVaOUhYQLCE2y4eWXUM4vbE/w2o1WKmldTf2V8E0VwtP
H1OVLrBZHfQjb7QCEtkSxPFBe9EBD5aIKBVUFBRAvAJvnUnBLwL5cJ3OqVFQ9JShIlTX86e1THPZ
WQ9D7iNOK0LsER1BjLccDideqjTme9rbdJ0r+k0eePBiEZA/9YBAQSm0EK5O1rxsUsMeWPGYvB5F
nWFoNH/KbWuHq2k7euI0go0o9uToLEgGZxcgMsh9LBIAEB8LCjK9bdeZXpbmvnPzspGRaBpGKpzf
dlgcgeRAV78kjF/WTSv0moYWNSO2r+u76efldIiCu7uWRs159PVtatptwlaRI65n63m6DYIs3q7/
2t3rqFYU/P8tDQq8mPFdSTZUrY1r5PGh2yUQFc8lwjmVGpOV4mjMuIH4AaMKCUFxCXYHQnrzPFd4
K8WjdF8ClOUB1aO3w2yjH0Xhe5r20LO4lxyLyQIJSd38Hd9b/uJdczVZnfNx7DdicgmdUUaOu4xa
CzJkkUXwt10PwQ5c3Tcb7wHyzUcWkzOthJcjnkiCiz904qZIIce2rX1B2UEX29bYcmJSqpiBhgxO
uJUNmlLiR01weEYXMEKSSMCSYxxEPsV+WpY7HtALcnx0yJx5LeSDQAeoylknkJCx4uOwgzehDKEr
ap0YMR2QZ35h24m0MOSbg8kcqDhoyC9Mc33bBUKS5xS1ev9DAItYHRU5ATGQid5Is3I26K7sOIxi
CP7/yzja/mdi5sr+4vj8yxfn6/ttHbes1/Ia2IsHgvDhDWlY+CVsyEtdPzONa7JRC8+UzMlN+55J
tupXCeiIRwOJf/l+J8bZDtYwvy2L9F5FGA8IHY2qvRoUUX9O1o1k3w56Jl2/3u916wgZA7+MZA//
RxNe6BPUqy5ersezSwEDwoX/FpDSZ/+ZmbSBEovaXovyozurOEPvZ+tWIRUmytwazMXaofboAnul
kfat/JMLIOCf3yss9SDvJvmzbSAdiDTv6MUfGvT1WAcb27yw6czbiEYzp/UnXcIpbTi5KgQ1GVbN
usn/pX37Jj2aHT3rVLPyEwCBYlrJgEzI5kD9d6RQUI0BsFMF36fPn5RW2BJojnVp+f/LOvOlhomq
usXV9d8Phs4iEsRTC7b5i990ha8brpth7bZyc1N++pxD56Ih5u5bNF6xltd16NHgAar9DS29NTLZ
C9izA1x0WD/P2H/5p3t5APiAJCI6ph2M8GPLZDvhVseHN2viN3FsjkXYh52xaX9kDWVilXvKCnBO
9WvGlCuvS0D6peDrUamkKznZgQmdjGCak5iJZez069zEKAZPaciPkbopWAT+jqnom4v4Toi00fPa
wobDT6p8hoLdpAItfGdvVkXRbFMTrqE0S7y8kDIedCKN2Y98e07CIZguzRCnF90/WGV+aC+azyi9
yQprC7CJh8Eoct/9dbw7yG4YczC0NAZRh9naaAZm8Pg3hLhOl6jel/+QRIfku69hy7tecIeRvWuI
Wf0HGPj/5c7AUUY7dRpyL/z1CvtlHWGKHDkxNesIPyZSFj8s71awMWl8TKxJBLVL6m3EtF1hCuDG
Q4Srd7fkVHodu0AjmsGobI/QvnSthn7iwQqpDLBchrI9bU81g8APFDZTpTPIHnBX6SbNB7oEPuRn
BlFlGAeMV3fqs+Vl13NH6DovOgOGLU2P+gXd0ScbhIosmxaGCXLwii97abtoNtW+kX/zGcNnsGpt
mIR0+qWj/EN1sHtaIsXjD3ZXRZznAoom8MIzjGu7AgZh7HjgZ9iYOuXX25ohtXJDOzrq4qbUQzoJ
/8QK6Q09COTxU4LYYL2uq3bxRsIaqgLauUc3xUCalDqngcyyeDIF3Pgqr3BJmgZb8iIe0cBjPAnz
2EqNGCkdHM99QwdY1N/xA6RTU1tvzoyVxDaWy2GnbVKaHzcwr+mgA2YrsqpSIPFsbccMTQuhvR2u
dnQaXXgU9BW51IMj6hP7Pfsj5/CFODXgpOeLKfDCurtR6Cl+md0dbaSAfCwe0dJg+s/2dFtzg3Og
1fXfHe40P2Q1mV0pXs78wlvzyoHuKSG3aUk20v+ItMyxqCWueY9AmtvkN4aQrzdsO6xmuGGnlHMQ
GuJNVLF81cwhha+Evr0kka9uBCwlx1oUd8aZ8sI62y9qhMb9zn5YQoWlEk8bMdUjTS6DoXjVA4Uw
NxLCrFJ2CPYqR26eoBbub+n0zlEtcMb4ht8MNwXxc7IkDuoULFEUUrWlsw5NHYXNjJLKa2fWxnOC
rbQBN+PVhaBtgT7Y3ulD8yZJq9lU176s2PYifEkibUWP4Vc9WiZZC5uVS2INTGPi/4Dc6f+ZoqhG
WOjE+tNH/S7m8AIHRvM5PRNK6iXb2s1pb6hvVj7ZqGwptomZi8Uln9PSg34sDdNg4Nw5oODssUpn
OUD57sSEitdVhMX7zyjx18doSN6RfNR0uHezwzzQWQK39F0VhhRfyfP+l+t2uQLD3BVAMmzzuUHs
sfpQlIngGuq1+lpn1sOEjZdypqgcCeNbCMnQioref5TLvXG/INc7mrYBtE5a4VetXkVIY/FtNsB4
G5i4Ijk1dEQQTycYu7RR7DtqyEO7oXDBp68awAIVwGjYATLHo1XTOXD9So9YhqGz/iLRVVSzM0Rd
baOQuBhvhUNOinZi0YJYU/ozAYYOXgSBIAHWu2zL8p47sCN6J38FdS56hury/E4SmVjD0iEKQII2
wLmIW3z9PSP/lJZDuXlrY+OS8U5+EGr2kC3lhjKR6z4kcpkK+m9gK3a3U0zBafmmw3VloAZ8tPbX
ci1LIF7un+ctPrBbXu/oCcqYPosQb160D+YSljiK1T4omd68Kjh8giHMXqEHBkoIuJPxI6kqIYp2
oBagHXVnaMo62piJgGF7ImX1h48+DK+NzEz9jiAQM1FCLrZMPJj73Ow/C/01fSG/oy/pn10oSFl+
6gu84YfyZfc0jLcIZq04ZecvjqYS4wjo051ANeCZYQyZeXvKuvxSjhU0Yv7wsQIaCxbjUxPu/W2u
z4/Nou6XrFONpEpRKP4kd6mHJfBpfILpIkKV8YhHopYYNLSa8BKRo/cP3zltNF22hbgtxAhlcDT6
qgmzuaLGky2UzBrPpRj5AAi9kpASCU+2iGH4ZgD7p+nf67pgOQiILlB4oSh4ihP1cfnveTEZoq7o
kwUn2c4ffH3wk8JaLNG+N7T2asYRhDMyty+avZGDpr+VPgcHT1EUd7o4di/LW/awnN3DQHCdKUYA
aBcYgyNQUNWVuU8T+nFoJ+tweOeQRKdZM8x/op2HmFjTcz5A2zuAFGIMHxmiEU82J+FYUjhr0u9Q
5Ci2c3tnFWeMHialher9xUQ54vOkiafoxa9D2TRZHJRtyj4u6u/Wpp3as4MHOd6BFaGKA/WpPynk
wTZY4ba1b02FPi/dcmRkzW5dzFQkYfU3+gBe3Pp9JlvJNTXBsdficp884gxYSHimJNrUzjDRxYkj
SG8e2aIIy4LzSKaX6eN3TUuA2gIT1awuRDsITOigsiVkAEb+dv/knrSItMa/KiHJi3rcRC8oYxLd
YZCnq6CaHIndZdaysX3D54jZzxraCAyehro1Eit3RC4IyBO4ozLj1D2lRrce++P3Heoswb851mNv
E70H9Q+5f7mWy2XAIG8kL9FDgExkNXtD/dnP0v1ko18lkeO4C52tVTQv9qIGM6X9gCJsHGbeaKls
/WSmK9oqTQpOhNHLPuSepYQSlQghEVDNNyTrtpt1Wb8Oc5+Zj/fba7X6crSjt9nTYb6MalANobPs
4zGxztETS9hT+BdfUKWgpKp3ZN6IflTF9E3Leql5yiRuatIc13i2t+fBvnQ/TmrB7EqN+nMhMYC0
DUzHqhXk3bVI64eSutYrrdQD3gZAjZ+N6CaqDzO/1WXSA9YsqQ+q+jmg+xxv/trtnjZLubkNLOS4
gZBcSj22pb+oSiKe/CXjTRAtpGj8GVnxQGFp8XuvMTgClPk1aWsXHPauJqJVKYbvV3jvb3QckN/Y
0N7z+jbKvmcQxem3dTuaAUgPgJE+SyVtv3M/mnk/xddIGwpYIyYjx6kfC+IMAiZwPlQNcoMZ9/hU
9ja3ykywjJS6P8bcqT4we1r2yy4qdYEGyrhJ4dQXH5ejpxQclm1jnj8PNvSbM7p9oFQ8uabPdWWa
jjacYzP2azCjDG3gMy3zWCH12xqpYbh09+z9jzdHuY6G8b+MlXqehE20a+0HqtmwoYiO1j5mVGpl
Q1Dh664Mp3jz5BmuJ8MbKEayjSYZeI0CZGiu2K1OzfxBvusNGzDVIzEdas3R+cPTVDGUY+lFOcoL
mBgWNhKNpCYG/tbOePD0rOk04+GbqUaRhoBNrl+8o/Z2lte4Ut7BUFTho9ZM2aN3pjJ3S2u4x4YR
bncyjnnMSg7oexRdn16wu7dI4wfob+C9HH6W4gu7Vra6b8+twUvsYfNLg8KHa5wvBdjLl2qkKffu
3VK/BLVWP9QP0sPqBi9nFdABkcb/6w5LVRswodt1+noo4xfVW72XObpqjmAtqvmMk671gndG6McE
kSmXbXh9LwTEpbqMgINyP3BdyjExQrj2M5Gnaph+FsQYdZnUwLzKL/mqcIP7yuoc8TOQuquqSmfX
1/zsPHF0QrEAlIr0fQ4FmKnClFtjoTHI6Vr/B+/9nmmo0sZet01imu3JeQG3wJEyrQ+wb6DUFGQz
bBYCVBUDhFUCih6qUg+QgoNFdZj6MF3F06gP428ufVWR/ocQEjcbIJsTqKN3yVyhlEA+0ZBunQnZ
TFU7Ac1wk4KHV1EZruGIKon0B4ee6TlbY40Ahq+pdTns1uoQ6xuWTZN4FXsciNxyKM4n4wCVuEKx
k0ZGAznjdpHvuY9p1bVZ+Ia3PrNv8OfTTUoBF5zolJ3k7cScBwHcmYlYDpON3nVIsCbE+19pngO7
Mh7op8iIxF7qOlC4Kmya8Eu2Ck2oqZWP7fmzfOlgD261LebqXcCD9PfVC+HulKz5vqtogoTIpYVc
KCgC/qE/+LIGvMFJK2eAZjTDgCElNJVUSKNfnfFVSMrOyfZcDtMD6yRPXjR1gQBlg7g66i+h1+/R
DF1h0gh1dXI8jknr1s/od1bQY1Bat6FRmXz2xrjxmGc983VQDNd94HtriI+lTkLHDhxkq4WYV77Z
O1/o0oHVn6gn0VoabIcefcgQKtm/hw6sB/c6PgsUwGJOj5k7iW+TYGHymCZL8gd62pys6HwwqgET
9pBPEhaV6moRfDmaykNt8thvT9dSgzv78HQmRDHm4+hIoMQs1arbqqONc4oLG04iR4dY5P4g8xeV
KKpMwRierv46+PG0cEcB5tB3NqtJPJ0LWP/Ia1/DUKl5UcKs35kSOKtRz/P3Lq9/H+lqzqQXQ4Vq
EvgsyRf7X7xHP1hpK7icxxA0y1eTUdbQAUkKD6IxEqPaN98Kin6/qxVwQorwbZN7FLfXPY6MCuUL
48BiSCT043KygTjppsW8kT8fHqAsNbB5xzpkfarEsEDh1EbLuaQraOMIfjRTiHsh5c9yCpPiWLGz
73BHeu1/oGeLASEZ1BYF+IOT5fxuMIUsWJTehmG1K6b8xJ/52Wlfpyx2Edq/xjlAMhP80XcsCHuq
YVq+ozdnIjSDj/97kCg79578L1UmfLRt5wFUDpoDYAStHWGvEqt5ANVfsy2Ie70JFJUExl9ShaMj
1i+FDJNKYvarVw0iVVPBzXU1yeyXS+WiDKm8VVbUvmiD4mtEUfRwA9++1OS+8p7TkhXvgDb8pbl7
MEgo43BfOPPOWyNQMiN9X9aZKvIjlemoNckHwGKKYBaECbygHSdS94i4GS5h4PKeGTD0y6leVxTZ
z4bsGJwI4ELxIw6rStKU/En3ZjbvGdgmvrA6dpjc6wMjV87l/If5m6VCeDoDUhoHCbQuu4AQMNwX
5Mcwnv1h8gx1egg7OGV8Uekhh3McQ0IO3BzqNHewAixuP0Ql/5wUHKOzj0V1i3JNVJqjcJ0oktsM
/iMsrcg7uQ4ze46eYas8j4qL96TaYfpbRa/cyH3gYhJvJjHcgRBYEMeU8a0JvJXHjvjjqm6IL3p5
sQSuU1N8fDJaaviF9Y/995m1TQERoiUoioZ4O0efEWh5AVed4j7DIV7gt5n7paqpL2wy4E144D1M
k/D29ZFr28zpPwmCAtVy95wPeF7NfHALZ6TVtdNepk897iaVdOZWIGSMSMRA9nl08RYyeamOux92
ZBvdtFG1z6k2HudBDK26BK9zKlFHmzqK25GGtPjTi1V6xw5+Rp4Rl/bGvmpMd5a1T4WvzpBProVM
gm4WYQF9XyOafrMm4RIkSrpEHHdHhq46IM2uDAOzHqqw6I9cIJKF0h9pYm/WzzXS5sk4oL/pTB8K
TpaRldr+hzkuMVzM6tfN2t2U5LNcQiH/6MLsMk/vUpyZZQOK3JGf8YP933VqJwnKEnS6ecMT0En6
SZYvpioMS28K+273jaYYnXWnjrgQL3IO2GxpiHAlLPeayCL0EdEm4J81c2Old4qcvhKu2IbWO+lp
QHbSe856iVjuBA04zySpcHtS+lWCyoFr+1P0CblZOlnkV0Gg3KgPuzOfMYxqmXKvworKTkW1EUZf
xbxgTTbk34pYuxUq+CUZoQTbKoLztd15jzg6/X1pOdg83gDpR16PEAhO6JbrOF+/aLHvIPjsESMX
LgXYvHFf6A+YCsHptzyyFwoUScFBhd4NqkaGqkvk1zb3r+YBVMhO6av3YdzWRgVTlwnIKgIHJVPR
2Z9cpMtsaCVDWrZwsjGckWncpMKskkLd9BpAzD/iE2j2XHFYztw5cUx8mvU47IY8aRz8x8KHhN2P
OIrOOwC210y2XvdBBictij6G7yhi+4G4WTYyx0U4SDQcOBJHvwJ+nPFFv5XY3tXyR9OEm/TeWoqL
XPVPgM5urU2/V0pcE5GblFBNIcXPUz+mO8sUI+cjCjqa3XnZOzKk/M+i6t3HPGSlx5e0/Y6Hlcb3
mEDdjZlpsscstPCCTEB3A4gMJ3QHtE1Om/ffAVdOrDt6iciy0zkzYeGSBSyFy1Ma+ZszMqEo+qJE
gklY3oLmmfdXx8TKybIiTFMP+tmFDshSf7+BP9/liIiR4lR4MIgmnF0LGqIE0eqjOTs/1LUHkRTh
7WNZ41PAWuDom7UuR76pjR8iaKpVfDmejWv/lj5qpnmOLDC00ubQRfR6+Rote9PF+DL0EMLUaUg4
KY9OJhyQTG2F/UZE0KiBGVkGBsM9AyS+FED/pOjDcG8ois1IYxJR0U8IVDFaXOYkfcZ/Wy9xEYk/
U7BQDvqibEX4WbaO35DtJ8kxyXOoXb3vcjgRew4O8eJDAUnoMA4Uq+cu4n0XJqXgBf9wpn0j/VD0
llFtUtUYX4klOeCUFh7nYT01Z7s1c9vlfn/A+1piN+w5x9P2c2VboPFRuSAwcQpLjgD14dhrFJVJ
J18ayD4ssoVwxQtgP16FYVPMMqId5hlMBa7DStIQWgySQPYoee1aiPXAc7RYEDmkvm+Zdbhjy5KP
5e6POqrTbuvY1H/QO5Op2YNWmHSRUWhw2hkIBJJc9OGwwyEZYBEtVZpvWteOX1kHKEEP0EPO8Sy5
GNesUIVN4bzczBrmZw8/gLTuqVO9UDHa15AZQYYyQPg+R3KVC950Fv89H3COpEicGqDnQn8YAGVu
TEMKXy7NfJyZynWRX27k6MbphslvFx93MDlEYrrZUv+cJNM8KdG8h/k+zUS419LAYw5fiY//i3C2
yR0faqbBMht7vwGfLvwRrvG/BmQke5VMo9NV7IENrt3KuSfuH0Qcx2/sP6CSbKUKqZFZlziWzuxI
zJvyForlsUpJZy6+KJ5Zn0f+IBGFBvjInAdfi8BnhMbSrTQFRvJ7eSxMYx1XPijo/9Giamw+ldcq
Udo5lZhgbV1dzVefGqBO4nAiSiMVMf9exvqjUarQIlxK7LbRoo3LuLwBx1x8pjgm+7+U/IrjMEFD
cAqnMly335eSMJ7bBSK7ziUEeDg+sDxxOxqoIzibpxRDvlimbZ3bzezQSWe5iUrh+e+ewY+H6s7m
u1eDu4lvlfsD+LAY1Y0J3I7oUbeKFqDSX/X5WatAB+TXpFq2YiB6aiM1yk2pyszddyYnTGFm6dQ0
nYnOn+pZePfOLjeCTqp2aH/zwc+QUafjp07q9+Z62k5ukNsG6/yAItKxf/bP1v1t7DjUWmAZZP4Z
W831xchbYxzWSEDDLt6fVkVY+2FBOBYwfxDpxpXsE/HkvqHHL4qTPdBSCr6FsebRc3tVcZqYPAsp
vgEqfvtw1lC9tDwYuGUbItMv42fcGb+wChrM3+W2P4loWFwRZKlW1Hn78BVKQOfxD3o/IaiMmVQD
rNV/4XUAIbvPXHrf62YKT6OJvv5CXRaQ4TAVwNHDeTgxf6NekYJdP9Oya6vPnhIl//b9zSQ7yPG3
lhEgMWEnjcfruj5Y80TKrMiV/FRnTSHNJop6CG4unvShN+lpK9qe9oW7knRow0VsKbnwgpHFuB65
BRuCe7YBjZoFB9MJl0Fsjwaps84kao6/p86ShH43qelsKSS8ft13A1U46GMtV4zcX9nl7LlEZ4FV
aosDxh46cGM6k8Nj+Aw13/XVC4azah7aEp6fGydQ3EERxYeiWONFCfrofi/3+pWfKIBj8K5DWnc4
EkdKeTW2DhVVjEJqfEpvTWA8bUcyDgRoY56nFJ01WSXNSzKY0dqMirWYxjGGrYuXn26NkzFxn1jd
5Zo0TfOcB49Ffs81qqUCYuwrHx8aW5AK13CQxO4tqk5wuk/XAuVZFXfq9rl2N+vPd0Y1Rtg7CnTq
cRBPiy/i/b6h1lkCJeRDZSYwUkiy8VS6KtBVpZCPs6La7fbNTu+1VVFGdzZggcE/Lr08sTbypdca
eVWWhtiTDU2yNZpGDaCZpex7cpH9wdQ6mU1bb2Q7f5DEwThPK9w/BzxwkBB/hVVt2QBMX4TLIyWX
aJp6ydQ+ZC1sann9Pz53kRg3YF5e8JBmNMSW14rREbFk+NRe68wg92tTka/SEFWwqSXSMCJj95vh
Zmr+MW2awpb+c9YqHMGtaixW/bGGxU2YnL3RLtAUjQfTTw2/mP6LPf3s5PnPMZV3z49JpLM7AbI1
9CznM5hHWLzG0Al+egxoTdVkrWZMMRwKgzQaDyXfPGS8+Jw8mMFLgVs39dfpA2tyzC9jdzDQvAfo
kPdjiHKWZkfPJLpl7h7o5VebWWMztcOH0OnrKA22x121YshWkjbz6kLd8SsRE7y6x9nVV3qohg/V
kte6Ai73X8+XPDJ8660TWqlzmS4tAaHxO+9LDxuvRvKnpnFgoeQXC3qCow5u+0tEXr5exGiBgnBv
8BxlIinzHlvfY4AYe2musCQnotU4jsP6oZTpmp3Sbs5WHpUXQ5NPOAy8nW5eH68O3ZrNrZiqokvL
kYn5pN+9OH214t+IMX3hmZ375ii3ArNjxL+rKK9uVpmDshB2ytJmoFyxa7/1rM4Amj9Zrkf+Wmk5
TikInc/P+AQIucxNkPWaSS3RE8bZ14lT7qJU0My1DopEaKMw7X95+7DTE1OoSbatpfq26D1qh0Ag
u7P68h/z+9mN2vH0LaMy5FhnseqkvDMEIeyfXBrgmbNJ/eevveDIZpP5xLWmdef/aRTD8TClVoM3
EhmTsU7xgrzCGyeNMzf/LhP/aUCHqUSNoSEVwMu97h5d1+j3xoil+0XlX/HpuwIjjalTBc4WRi25
tUqsfxI112jDgKLdQ80gojIAnBV2jrpcVDxvaV4zRH1XtTDBARvB3u28vPr2bb3HgJvXeeWYabSU
MaguqvwLZsWKw6F3yVD+glQuhW+la3K3TG0NVDztC1xXRmCHznWiB2LAuu8ebeb58dhpC0onlm7K
uqthKr4wVvBwnyBxb86QR6ugN+ig2fVqTUfHMN+6j6xFUl++MK5Yb3Eb3PMJNGUK/7srXl3gN5BM
aIC4TUCixbnuXCDsifKYHFts4LuChOn3BWodxLoE3sReD/372XJCdb9g5LsfdNqD+pFicv25tBu5
729A/+3wJ93ScRS1ugOma9Co+Y6XUHxIeA4IWad8TcroHpP460X524s24WkudZDH3JnRf6IHNPjc
oIWWSYVzM9f/E8oP7Woqxm7EAn//e1A19LfFsJaiUsTfo1iQK0eHD5daNIgyrd0gK3FuIlp0zVAN
nzX2bG78Bg5yuuGnqOnQI119QAjgiOZY+ofFWbEaI5gOZ6pXl6VZbz4rXK995rJDTJAEGRP5YaF/
oeLsUUIZ8SApn9jcpJp9qbn0oRmQxie4coN7SY0q8XirGotstUe8jC9KH+b1xiqt60ok8cqeecKq
OU1DvS5PEvrwVk3gc1MzvntiwbRwAn8r2ok6nXDNUOGv2zdAXHTTTAUSNUDO4zJefpI27sFQbikU
kgLPTk1XZFGlS7HMmjY0nTSsnz2NUfyTyJVskAXzX+uOqwMd+jOtnrLx8mBCQHLbr8+1KPJSw31A
iuejqaDj6hENcaa8XQQZMT20p5uoYu/9ivgRXdVDJVIfaxNOsiZL1Oi9Ujhgq6FuDKI3titV+6R7
CXFjVYrQRGKDI7sA/v0/9S4LBCZ8eXljcef3aiowMTX0DYrOHdRtgEYBo1FKEqAxjpaf7IKGDDYJ
ypLGwqYWlh8OEQBdqDSUhlbKJrND7gIIDOdCSiuKIJXQEpg4rw3mF9YpezV0ddiJoGfczIveQsEU
7wR8YYEmiQjCExVE4saZIQHmSX0glGFJzBatyos8tepRQ4UjC1j/cH0PrcJ7eQLKiWBMff34zO7C
LEMxzRUzCvXCg7DLkUw24mcFz+JzP5862ehA9JKrmnP6yPmVO5ypwKBKwMGj+PQ0X9N1LiVIdbVX
5XkV0F/fVcRbM5abig2AtKmY7xz0J0rB9NDdMIRdFAwC12UGaLb/OzcSv5jyHdwPIzXLxi5puwmw
WUFSzYaREPlDE9/qkWx+53JZe+XrAvLuuqiAxrcWp8WMQVfJr+aeRHQZ5E8QlLR/6UeJDq0zsqDm
x13Cp+4YD+TT/yQIUNzRX0fXLKgPi5zr0xnSehrePsXrh5Eg6Gxp/Ze4XpS787mqWtImJu/AIyio
+9M86+Ye3IBEMhVUUjdjfaNh89sJh50jiGGP/45lJXphS+eOM0SgZo8BltkgGObC5Z45NYmEqAaL
jXOUovrY3m1+pnO+B0RJKmsm5Qa245erA7fpoAcwSLJ5CjM7YxpOwd/UV+i1E8yWsGBkUHE0ritl
K91wWBpzZXCzRxp+0w432u1WJU4l0px/jI4hHdzx+cgzoO2LqsI0yrRee0dF2g0ea5UlDFs31BKV
cEFtqWfVpUxRsuTY5dTnEO+rtFGRtD7riyBM195iQWpc7J36q2dt7Rpp7sVhjVjWL2b+l/jglV3E
wMzOByYciQvLOKa3kgRuYeYkHdvaOZxCmUNtIhvtqCm3kWOlIPCoZltJFg1BdBhO+qnCOYZwpaoD
1ycqHvfFGE76Od8Hh6yTrO3pp7AVzr8hEMg/ZRPoS0rtXuFhdQSZj/r+zsrAeebsyoTmqqTb1Z8N
Jbsm+oHsmfePMDWt6KDoXG4NoMRRoAZhrt3PhRTmUMGPgDcEti3NInuoIfqKRiHyoRNK3kmiNOU0
/yE9oEVxR16PnfPrER3SiPOkMW0Trp8MIt91xMuDexoMi8H3PMDktLP/qa00orWD8kruf+euMbq+
jLeEbeymGyTU/eO18DfHUoJwSbvjl65gei7ift0Y8lQ5EA/CNhFrlk8EDHZBVOdQtlI1wV0os5qk
FNtX0ZR8ROOBoBlm0gLoWQAZ5cofr8oFLXGlrOzieo0YAI2oYlhnuvUlZm3HxmTVhLwfNMHp7jF+
hh1jyQMz2fqSvqEmN7cdCSSlNnJUUee58HqiyPLh3LNX9319+/2fCmJX4lCR0sCbPzx220J/lIuU
lOIaTz99Aj4gPG8Jlp+6qz77VsFCm9W50L3u8j838bl40E7k6Qox4UKlz9XzUCT3IqgF9usP7NHy
+jF7R3koH80bzrHo0yYu9GQBAwm9iEE2Y1RovityfaDYTZLyty4Q18k+YVmV5xJQGKvBKHEj0g7K
DjjLXdVc2oMgD7kGlpvK8+hg1FMsGI7sVKSzW0PBbqBhA2yV+2VKEiniPRvtVb30IYe2ZfrkgWvv
ofaAXluj1N53HeflMvoc6/yc2h5E493HL5Tz6tuZvCCypRIIddWFDAQDfHqpad69TLc+o+Y1nJCL
2aaPVgx62FMGu85HdNS9vdMYNB9tx+r3Ij7HSkdfkYlYY6oIGXir4GlY68aXUK2uo5uZ2ZSViZSZ
ePLgtc1S/sZ6ODdouHf6hWyG6wYXtUoaWypgNEYnY2PlNEHCLhRE2QfqPquD86hRMBFKXs9gUwgJ
zRBZVgX6u/UGqs8SfecqDYISgbf7oQdVPcMmGM+2kg/sQTN+r50vVQ86yykSB4R6Y4gFLAj5lhJQ
o36i22kEo32I//jEq+2VKEiR7sHnwfTH96Ee6wt0jdtS0sq1YF6jCZzTeA4COeUb9K6eIMIVq6bK
Y0f9/gK1CaTL1NKOIfeQsYTDYjaOPkBcwOG176gLboIOydNzpZ+VeOPXNFrJp9AFvxE7qSblyjvD
DQYsuKlfabiuC1pe5BF2/tBXSoQ18KPB69X57cU2QJ8rZwrZwR2fELZOsU+/vITJaCG/yRB0l26x
wBciEfy3CwKY6AFslCNxVsYgD4Z+zgLAydHAuNlYvknVOjgcpWm8fYh6WaQr+PugEDfwwfXqX4Bo
OdGqvojf/KBZaOVXlhE47X8VKK1wAfWtQLCg2wSO2dXlKD+otvjZePlWLkciINXrJuJbDzUUtq5B
aLfIuZUYXKUefA1YwQtpYxW1lSYbRD9Zirs9RAltKY7ughk7JhM1Gd20xesJz//VWus/eXB6Wqk8
NHfXlHf2ID+QD6gA9uEtiLgH+T9kvUThO9+M9XfOi2XgvAKN4yq54j1Ocz3A2+YZVtT3CUUUAF17
Sv2hmhuTDa5/oV62G6U3pafuk05uNTTs/v81vUgEZ0zFYIHZxrwnN2m38WnWVPMg1zJKt8GTkc6w
i6AmyMPfVhnrjpcf6TwNS9o/0DLu58XphVc7PlWMNWny2OG6dCMQ+Ujbww0fGVJLdcbzIYRo7grj
p+BganHAMb+wK1pYETMAQOv3Hbr8ChfKQevnLmrplwy4Gb5UnRjzZrD9vJn3A2GvVGn1d8lfWRZe
bpJ+ZIDZHbF2RqacY7M1ZscqTO7HJ5YfVwUQbhyavSAfNby+FSsF5aH0SWjFQa/IpWn0qtllt+s1
Mvs5gJJzFwrNuBMv6fuyQRhrFu9q/0YU2vc1faI1Ucey7vdUysrLJyBbCp2eVrmUou4YFBzHzoNl
HL0o/68LhfkLgQ4h79+3cl3ExnMW63f8V8ivjDyZUdsfWagjbz2hnHCKKxZFBG1cRkP8gv024ROh
b8BcEv4EXK1ftml0a2HKGBy4aIJFVRAwazkkSAVMfZd0OTVmPItqH9pbFWhStruCB4Y6BraznI2T
eKM6UL7HtL443yyWZn+UeuhuIi2U4bX59gB4bGmx3AtC4JrVm26wTzXDxh5rsNunIgXnn0MY3CUO
IX2Enzk/Wns4d71Du9gCS5GutSYqeqiAXnJ8p6REPy56DeTIsS5WHSwdNTUSlK8LdgAnwpQLWRYn
ETZuwdnE91obmVhPvXjpTRuTkrJItk738IjTdNjVzCPCsnxEfz49Hwju9NKBx/V9AlEXYwHzJZ2W
uQ0tfKT5eKevrxfpZUvNqS4NCWrrUKP4pDvObHwOARNc1lBu97Ecal1uwXdLRX1vebXqDBbhKuU5
MqZ3RUZnlP5Aj3VAnDdlmXMzrMwrgm9aAVPot96N9oH6s5rLbPls73szx322j3bouS/Dgf1sH/zd
yzavrBuAMomKIGRZNg84Ijhyl3407dyg6/ZdwBHGkYXVzZpnbEYD+j0O1Nz9n5cXUCOKEPOOpHpT
2xWdN1KxCg6c+Q71GO4pWRJMWzkG/6vff0LwcydIVu9iZxtODm1yojxpQGSDexQQ1mieTjCjYuOX
tc7EsAPg3Y+kLF65IhwW9vkQQMqKnoKcB/0pxGNtFerDWgAZYa9CAnzpG3ksZL1dpvkttCJR/oy5
SL+p+GtlYczAd25J01xNJWege+/dOwKWHdtc7hBak4BkNnJrcmSqxIPChCCNCZWaoMy17vHkkTv6
ifRUvHodZ1JWXx4hphS8rJkCTAWX0jt+RtyKgPbXvb+NSfxbeoftIxrp+oXshg1d2eNB3Hx/hvSV
f58L8f8De+13bMLeY0Q2Je5rwt4CJCo9uV01b3Z6tjJ3yDTTkmoUHBlqDO9lc1RwTiCy5THEmALa
V13RCV+dzQhq+Wc9Gwg61jcbYmda7o2MdIoknoEOAur8plD5ccdafSXbUO3+KwpNdGgegRryIHrW
Fz/CPFMKC05c40TayYnjPgJ6v2YAMDxkYHGoO2bf0dSAt5pfmbtifBeS0+iaHAG0ZZOqXfiaq7Uq
FkYbhXjBV0WdLRi0DojjrpfOrM+le/rPNq0EU80REAGHPVZqDnOsTayS6pfUIfjdid0iBYnm1/ep
tsaZO1eQGyBxyizZhbip7FBtN5i96itMSPDftyEq43Xgn3q/fDd6PTHQXP6YOgRZjaLfK0Tvaa/t
bNy+13CiKd6Em6LpjuvLeasyEYZzpV2nmcA87vyfx7QC2RAL6CEipGcaLqRc/6vmJ7XRF3fx1zha
QotzphI9lZHkMiaJbTE+n7+qrrerpdwuvwgb62gQXYn7G7ATq/GIFPngH/go3zmRQhCL4nFwOIFK
QWqqdZQLTUsPS6xOP2lZvSig8Ic4IWGbioRY8GQqQiTzI2FQgP0B47oDwatkixWfVYdhPaKWsczd
Z+lFBjIkOxKWIFJdLcHvrsNHhLI4DzEcyKJ5sgmz8yhSXlB7LUj05ORUzzu4JI7nP5S7/Krb+MxQ
Aj9ob5o8IQ+/1VYorscTM1qOWFBIOLwNUuG2sy+3MZ8/mOYaSH4GdSmiha9HsB+gKXE04n+oxuPP
n8rgnWhNXKIb1KW+ilMq/uieEOSbS6jJU+dPX41oQoKzrxE/tmiR8ebQGdd2vhAS+BNJT5xA3ZG1
dTFum22Y9NFYypfCMJdPjkcWN5z6FbjPEfSKWQF+a8YlZSy2VToc5B4az9ygbpuS23jrDNuAmSlp
Gm782NtN/8tvN7sYFsBB5AFUkiRi/FkxRZajTX+nOO6gDkRkuJl6JRVFqdFA3MKBZxjECkN3qtof
lsG+zXpYlVN46tyNHVtPLvyA+kuTbpYDkrcq3Zv8hoJ3WuQkf6sZaC+uMCITogXGt82QQJH8L9Jp
soboZJcq6b7DLlBBPlXL5jkmnbrAEIBiltzm8JuDtmGs3fPIFe7wgYoZqNiaPKnaGTVivzfYwgWU
Db8GZi/Yt39yW5qY+ZkSsSlJEccP9iSf06elBUP1NS4dxU/TK09jLOSziB11BKppOaytjwPNClDQ
li8mFSVCl8SwwLO7oqmRdRLkD678H7K1e/Bd61kYnMIUeZkE8qpx49H4uirDfncJ8c8p9bxWcZOK
Wk2XBVlpVUz8yw3o4w3baBqxi/gGxbJhXO1bSEPF7LGFisLg3ES+MHe6U2oCD2101VnyePkHhFxS
a4loioWxjTvnWdyUurLSw/f1Aj7j35bH6iUVT3UBukOAkrXKPZraZaE4itwzYpZsEDKYExkYLGn2
MM1bsmGXvidM68um0tszi+OVQiPAAKAkft0SD8oUsqK3SodN4S53x1XG31wEF52cNGOp8PVGaWSx
dBN13uo57HlUB1S3uCu9L6bCk4EK3zRYl58n9gvJeo873V7mvNPiIriq4r5iX+iqbWiDYGnhG90g
tTnMEVKr3ykwJgQM5JR5BKIW3Rc8aNgAL696UT7J5/qWhhtGCOYFYNzbHl/nz9uooULm7LWH6Wom
3lUTRFrzNHD0zOU66H6ENfiFaCLrL2qyd/lDHxxnDxRgrQudQfWJm78csBoUqfJ93wMIGm7kPMwG
+/nHFjpu31lpO0DT4VBU4j7br2Vd79VuGwdafI1SDtrFLgqQyuAS8rNu/D5sFUHkuqtb3+t4+OCy
EIjPjxOakaYZhpv/SEFg7nlYMwtbYd7vkO+Jtd2ZJY5wwUowzejs7t53Un4GTvDdc6eP+h0CFwgb
DsBqZDQ4CFdVTvpy7hXhj881CihJyyz5XgkfLjM8LuO4EaCZtRkL2ZUS95GDiSBHvZ6q9NZka2Pm
QFTKj9q97w20C8HpEs8oMb+7QXx14hXrJKoK488pv1K0jSHx/1QSOs553qr5wh+Tx0Eq1b7FPNIb
t7binnfnNzyKH/RmTLRLrbqDDhT9jDCQTbj1LO4aZT3zDA1iiuaszzJAieoI/SS17yEKhwvFjv1I
Yp2YeRSygVRqiYAvqZD+QfclOg4ogzEf3vPlYpfK3vZ3xpk/S5LihilDtjw2Acy9ytBfb5Rhtr9D
5896EYuT1Jk2dOdYv7tVlFnRAc2XDV7zdJdvSd6PorjpYrD9KpYW4L0yKMbjxOcIIiJgaIVN8JoW
RkRCSgb5KBnDj/pBpDbX9pe6I9mD72NNw9vPgR/wel/JcLzDhKkDVuDfGJy1CcQCprI0HyKQLD4I
WROWsctB4fik35meG1ur0LY5VIFjQsWYNqoXy8q6YOba/11g6VMcdxeAhFa5gE90MjMQQlq/AOm+
dAJqmiT1BNJsFvVVzeX34MaSkYUiq3OKc6EIiyy2VCTyNcG/+VynH9w6DRMo4INmjDa+W7UTMZ2Q
SEWIZcKQF5VkubpfXRhxf1R/ip3tplOY4u1c+idtpfSWFE5ODfHbisrCDw9YKy3z73eOD4jH0RCw
SCTe6Awb+/y9hjQklcBhjseCrGlDGEY9wweQYEXlX6SFTN4m7E41wRKFg6P7/RebHXZo48f6sMVK
Qs3ZVF9iRQDH7HDbUhMj1qIfVou9plpGQ/x8oPB6W6909LXwAPtUQaicuwOUU194wbnXhKwciBQz
ar80p2KNS7yMSG2Wlqg4ySEWh5tFlUNoVgiYZ582WS3v0W94eYWIbYQfID/ew313HDoXz4K7+v4i
KFph9n5Cqtjp4oFdLxwYEtDURYoVEEWtHp7oUJAhaSQ/7ZrfIjcN4uuy24n4Q6aeKgU/LtAgvMLt
j/kU4nMRT+8LK9BoFJTN9jwS4H3qmLf/+LkvQUAip0pggYs4Y4wj0wljbpbKE3XNfrqaD55Tw5r5
SIMmHmDeGceeIwYACLv4lUOJpo3I+3zna1LY/vvC62UKvRrQIJTUCF+vRuhwYfSeBdhyyBkN7lfz
f71AJeP9r1dDh/DCpqfbJp/hZNY7f6pLBKGc+6UsB4QR2Ev/HtY3Y3EE0XZlx0Mc92T8/ygGg1ry
A8HVCyF5dI0PfkoZZMxx7mNZTt2APkyDVf6QO+VpUnbDQAaT4J9TaHRfF58BU/1Y/rGb/BUKsWO6
9qjxdta502k6RzS9JtqdZbyfaj7Z3wVMZpCZhCNsZNfTbqxeG2+G41b4NC9kpeIzjyFupaFbqZaM
i4SzBRffPcDgUABYHMcaM6HwFZwWRkt81wWbIufFW8yQ/tLGyOPCNB87JZdJvDTd0vOI26z5V9HL
H+2cGVziRt6NdwlabAX521chepYccdIKgUfR0DhCp5W2pONJmXwf+jjcPwNzwY5K9RB91KFmWS2h
CCl5BIayZEba2bBQRR1+ENkNY7fPxQmTDwtmjkGZUmHBThpK32T2EyNicxJHxt1dOumCLN9TODil
Mzul/UkHaL7zD2wc0M566ys7M0XiOL+ei1v8q1Xp1kuQMlThnrNmNmKY7y3B7gc+QkDsv4p/Ivvz
QdXvREIUczud9PqkVvnCq89VA9tXDc2wsZmBVOR1CL1FVIjudqNWc4Awr3SwN/DuzoGepPJxflKZ
0G+6hJ3PUrMmJyK3J6B++USkAxOdR29LYw7kfP21r5K92qzACeOh3V42+BUSCkFs5vqONzXf0Gcl
Hb5spJxzsZnhtSXJ0hk3WwuJEH6Z3qmrz6m3w774XRDtloGVnjR/s+/r5BOeDaSIACHPtGhAEty8
zDuXxFCyP0N0lb94N/iomR1Ek+R+VlIC4NUGkBuoE4dViM1vwzn9c8a1IVbNa4u6jMjmM7qumZly
XPTxDr+5DkS1zf09LMO+X8pqdwCYvn9rQL8tCD2zALGEQOs3Hj74jucruR+gI6OunTDgmmNBJtt4
QA9bjex6j8S+aYuAOueGo+e+0w0e7Hgn2vL+vLQMW8n9tbvgSuy4vYvL3uk+4QnvmM2/asAOyCNM
qRqDcrUT6+YFLjduQ0/Q470sTScqVPQ/ZRTer/vvF3fuqT8OkSgNrS487v6ln6WrCP7ApOXMHmql
M0Ww8SexRIu/y+06+5n5MpwIRQC8RX9czbgq7Ojm2LDrecIXRGFUXsnxxS/sFSrxe683ucHjPW/I
+xdYQAly2UY7uN1i2iKchkaNwkO35dWF9L5KUQqLhST8xuIcGng45Fd8+Biga8zT64gFmQI5XyuM
L7O+0SZSEVr04N2RUh8+GwNhcdnHmxfeYHGZDCX1HMYdduugbhlbWcII5KpK8kQoyUvBPivM23px
JlQEK2zvavtPOylbgG1p6HaCYhdc3O/I8TFLAEOU1Z1CbIFg5JNxXfwe5Mzas8kVwu24RZ+OvZPP
4Ig1HpoygMsoZ4lBr6mTeeCRQs67RNsxxDBustA7J2lCiBOSKMXVpovsgxHoe7oMjj3IoEn/Z2yL
vaCgc9R1ot6u1RVOR4I00cSiHPFeSjvzfvJGV1HZbB2jyiomcmwgCId3OqY/mUHTboYDNSInCjuM
IrP7F+BTMjVTrKih8XaAzZbmAmtoZ9p9bsLxrL0DnSLRjOymX3l3lxB5Abp/sF/QzPVhG1qp4LAH
z5InPNYGwaDUc8++nSTMJujqH6QOmL9If6pdXVVQllaYrr5bA6P3LXBXR2MdPsJWTuVTZ/Y+chA/
58zV1flWyfK+3cKRUIKwcQeWpx/IDfYaJuvkJCc2368ci76derXvtfB6JwRMXfOKfHdyMa3pOw7o
b5MVY0psJwm3iqIqSDmpG2EzQEg0nFfDsCXPN4M7ffumB45os2JAg2jq4+ksrdLCwEJkR1z63p1N
WufAzBDWBTe8JrBRHIeH0UYiR5luZFBprz+zsB6qyHaCJanQa/Bf8oVYoLlKTL9FD4wgm/My3+yg
V+505STEq5+72o19dl/oakB+tZg7e+O0oUAnRFlqWstfZOJeSlVgGZYaXLLRKa5PtaYi+hgb4yoE
QUoZeZ9N6wkdDdLoFE9lNLma1JgOlh1iK1dVidsmNMZJF7mZN37TO49W4co4qamDh5GDABn9nRqz
i78ngLTtaBuzsBMx3FpE86g0N6D3llwSapUq7wqMVDW6LzkVpFxa45t14r+PyHNYR6hxwqkWCAR2
5cQtatqJWeJ9iB0+FTOz2p23ZWylZAiUArh+VlMa5Y87MqsEGcolLJ4+DnPLmwRnG3nQsJ44XiIG
TI9IHsjFaQhVaZ50gDIhbzxZtNreNKYVHPL0TPO9UW/hXSzlPVRsmgFzoTPs0z7jsoieKCZfpl6i
HZfbNEbOTiYawCYRlPlCdAvnDGxaCL/yTdLwte8CabBKrV0h6iNCL30MX5QpOFOKofA24NfJkIpO
+L1cUnb6NR70IlmncIl9VvJJvVy2H/wgqSG/wjw+Q6EqsgGvrz/WX/g1xnTVeML8zp/HdmpSHAFs
cUmos3Atp9LKBiYdKkr5y7ORw/g/ueTmc9xS9RjDlBeF+uBto68cd/lurzRWaGdbqxNJIw33Az0R
+QkULQv6sou/QC5Pd7/ux1m8tmOYhz08pzAZ52MvhlJ0ZzxTSqJ+OClqgAnQtbEMhaE0g5trEI0o
C4fAsekFmRf1tU2PrgV8JK5yc/KSevP0vmv1OyVPBMG9ASccaki28BCZGI7pJOWJ0KwB3DzNbNJb
nGL88GOGVJZqtFkoeI1ygqS5LmI+gDUPTQpeHH4wb9z+XstB1z+e10QkFbdb2Zn3aajNbQddiAvs
2U5wUNG/JXnroh0k2hHGTVdHZxq4KkgH30Zsjru1p5MZAmkqLQ7sj2uSr0ZrxeP22ARe5sQvE5Lh
b186Q/UyBzN9y4wrm6fn5ifuULW3SL555XR6RjCZ01/RyjAWbKl8MHdvnx/Y8OqBav7x3gb2RpW9
7u5f9qpU2xLc6e8O6hj0gfZXkN6orDpX/tUoGDvh/gGNG2sRYFlGxKIwwgHRQ/VlidHRzxMoK5OF
vEuYH5yKTflqGeWHmg4ySWpBt2FaDB8WFca04Rmd55jpdY0Qe1L2HYw8jFeOa/4F5SspWOFxJ9zA
Bh4wAotlBnj5CnnuLmnqfcsO+HgqsLl5YwOu0f4P7FKm2t09X8olLuPk3eYZu1Oj23KJLHQ8hyYF
xAod+EyMt66rTKIuScBFSgSoF0RV0GWHINUYpopYSH5juGcAfoQnFmlLsRal5Dh6ngKDVVSSKhpO
+XroGx5fwUqVl/BAWCctUwxGtR62zdpjuHZHdcUz3luMO4K+V/lSlnlv4NKKvswfuKPGkIEwPkoj
OapaiCVAdNz9b/eZ+HlUKIouuinv9Q6mMfL7GmsPQ833P1rkkCGrRvNP21bBmq25GbyAGsc+nGfu
Ny6ZjSKEEgxfPlez7QfoH5h51q9rzfvb951zYH5wM0tw2zE+mI3eO6MEQyJrPUQvo07wlI3Ed6Hj
FBdrZVrTmFPwVEbXYYzz4JcMaYNr8AyAJIHSEYvrr558OfGzfOzisNRQ+SiJj6PmuxtW9Ozi5Tu5
0gKZTTS2DAjqvesG2m5oY1kHRpgNydt3WpvZB72Nq6iDxgR8iHYsB4VGD5FISmgs2ZW4PYlxno4q
HzA+ez2lnUf3ghrIeiMOl6md5MFuzQrlIHjmD7SIOqaboJG2qBlNyt/x6vIMML1J6z3Cd9XAjNO6
fpc/6g7Frb6vBKnm1k4FoDWmPl8nzpm40qyYcrr3hKx2niYgzy8RAdSwJBM7TFBcJXbExQ6/1c8Z
JPGK16hf2q5mXCj/eCNfP2Fu9gBxrojAmpviUI+3B0ZOjL+RYS+XBqOwuU2ZKq5euj+LzLl4DMb8
AxHNkQlBDW1K7vEEVUiTUy+5tVew+6tgHVCTd0V6ixc+4ggt+I9D3hUhOlmWKRczhMqtf2HiB0uU
VYBBevJ6kwNw8SaJoPkFYV4aeL6bS6rkwWKpc8OA69kdeFqaSPQYAw4SMZuzngqoLm7zhq2xiDx4
HjP46XG7P/NfzxglH/tNq4mZp7fZu4RBOl7ERbYjPkmIszFm2ny1nCv6Zj0rgEk6wzYRTxd5xs06
xoY6H6oNg5gubRJ0XGma7D1e0K82PKoskvheVYOj36aA59SR9CU0La+Txaqdka8khGH0ZO8UAGLf
Gp4iLbOPigHoNOlof0gEB8StSUC3n+jMQ2gwTIQAC+mx/XS9lpDwykl7rpXhGovhHFTiEhSWy561
58svfQXVQdRxQ+SvFRY95LntKxZE6jC4dz8v+Jmw2WQjLLFa6XlIGABijHENrebRDqNdqpRPCZDf
GCEj364z+Y0S7TkIsjJVly5Q5m79WpfyMCWNPaESKrmEyy24oBk54Q+/EJTImw0a9uIvK/oGgv8o
vbDpngZe1eCoU51spnGb2wWIrdhXx5bh28KqRj03MhunNdoRKqjwJgBSFYmMjBWkxfjQd2MPyC9F
CXu37sjFnFPsikdiL2z5vzadn2aPxpqigw/cIm9LRVr7gcwi0AfoBCdQKzjcpuOcTdX19mlo3FvM
s6MLRme6vZOuPSFt68FZkzORb2i9qkQKF97radEaxaINrcVAoEPoPUY1o1adcFcb3qFrn+cGU3XV
XpRwyAQ68kn82n81DT06mPUdCXuAMWm4ti+CAwVVaILtTte7NmPU3RTipEOrcaDVT/QX+nCNFv1q
nDCHzLfjgu4bYplLp/vGQWFGkUyrzcptlTHoJ0HpaPfNW7nQ+9ryFb2VFaMEzOVvozw1+t5tsp7r
jYCHCrIMJqcgZ/7DUm1unF2fG6dZimWF/t4FB8cfZ9LTB/6x784dEmagnonCplviDuTJJbA8dNt+
njbbc1Iy9rxA0xvt9lVxbPPF7/R1/RFTlQeIj8bxeFS2IrWIt+7EuNT2LVOIdv/X1CwmJYehzoqL
F+cY+CpnFkOxCNHLxUZ0N7qJX+ntnSLDtchIrZpF8cpFTT8akVob56rvAEBwVFqHafvqsrb/bl1Z
aFJg3ntiG5eUDbs8nS7TvxuhJiNl+eykzfT+Tbiyoh2vttlrea8uUuzElCTosJPWYvAePQtWkSzS
GA9d6A6gPprayFUGGuPqJmrY9BfQv952+OJywS/I1BDVvR0QtCy9aBUycD48dbsQizKfbks5rhWd
6+uN1f4/m9TXT3KBkXHD/gEE/xOFSsQnwK2StAhoRlJ9OI7XCxwR26vnhMgPRUWge02tKx4B3cv0
kVclnGIT+gws55eSdq4/IDrD0bB91uZYCFC3Ype6Nn5bgHKgg8+Te3J03QuTC/8saaj7ryK1KSF3
s4ZH2PCTUhTQGJus43hUTHTBPuZVSEFMsQB5kHGwPCjH/C5HS4qgBYcrW8q/LlZ796zSafzAfc9/
MB5fCHBPEdG4kUgVOjgIXu5cpviCtebUp3ahnWPgvMkyLWlR5GSuU5bv0L/cVnSmiiDdW3uaDhSI
ElBDdag5jKJccAReSaimZP5lIYRV5lKcfYsNI509JQC1NI2+iVTus1X8CCm8vRMH9FcULGHnus+T
qHdQnNRODwCVWD0YvJVCZYa9VY3A2A8BtOfmKSoxEstBQyzoPVR+c+U6gvjQ3MfOEk5EPSrs1Nht
eYLappLHYCtFkatmertVSxx7NadQjMExGBiNOpOa/nGhelV5pqeHbufgdw90aPtxcz5vwsylWkvu
gMS0I4KyrAD8EMafqj4ZX5OHR5Y1286q6WK5zPYDqlilBH4EdnyE9VxYnzvjAOSZxhE2iFf1NLEG
LE8vWk8znF/CD7oC/U/X35ZfyWsXy3Ub5g7jE1rtcbvPLp96EBbSdbGP4qQQOo+auyKl2UWDXFIr
PlaegJ45WuR4VUWRNt7Z+YD2ZRUdCJ57ECwhzic9F32yD03B/0OYyrCm1h1UE7exUILmFj7qPKG7
mE35kMZopt7MfxSPEglfwyCjwN7er/ZWdway+2eQtjt7n7KrgRoEKZATiXq4CrRMrpfvpnvTVdhO
ipOxmyXmDUWB2zBFO73SW5HPmoO+2uVEbJdbReExOQSHgGuT72eyrmngtldMcBbpY8KSRR6ziesN
7gA2L0IYcS8nMUjPClBXnC4bkdJL/7uSEUQDT0ocd6NykvHnX6O0dN6Uujyx5ZT/aaJWTVzF7TLo
uPCwN03me16cNZuNMjdARH+rGxsiNZJ90Cwrff5qLs/XLK6IdQcWzv/Kr8K8lHii1MolAAOC2oPB
VL997Cv8VM4PWjOihTAsEUTdjMq0qHa5ovisZEktSYqdgQbBZLfYmF2ZziKEJKvamsUMjRr5oET1
2N3FU2kbsQHR8+mRKiS37OyPhHpD0xMvWqehAUIXpZZqpcx2y4CG8LbFRM+9U0R56qMWYMxEmsnC
EpiefG0Yn8i0mdn16oH30cbbAe4Rx4WeMN+pJJzdJNFX5YQ3J4R4R4t1jehKHetCRhu0De51mwfN
5PrZLKkUHMSnKHg4SFimWydlywuPenDIqBm9eDPQcWB/v/j5OxlkH+8DJSppU4EmKBl3x1j/AUCq
tbcNY4PQYCrKmLInqtJSEnwPUECxnfB8wVzCotAfmELNh+yxrmZ9vZ+qs5HPHNmOGS8nksxxNsVv
xo1uKEhXWPZWvckakzBAlHslsIHEOs7u6b8H1SQXp/pKGDWJ0DTgAk/GNKAVOUkt3IhZmrGJFlGv
PfWdg8usu/rR9/MxHZsyqW8DzlsfZHURV40ahY5KZ9dbK2oyDJN0AJC0xOeuRDoUsGMPJSGuWj57
9BnFUB6flhiKMr6RVtW/A/NB63/cx/2vxCt09/8e0rIvRdKZdx2qYDQb3n0fWGGD4NVIZY+E/Klm
QT0pBUanNkt0uLSG3q+s7P0l/igjcNGi76XZK0VVwTw47t37RuNmtu35M/R8dTAe3ktb1x5dAqZD
fhdSzF2+1vUe90ybutlavRfUkrdW1HCXvmBMkTYZQjvj1xZHL0pT7BIYtI5xjTDTu7VoeMIRv0Gi
ckiaLL+V4d1Pom2Vtb/TcLfwqCCSFVe57grObR1P6va2N9BPNaH0wsXtvYBQcOQHOYZA/LdTg6SH
JHpJXYcHA5Ive7XAwG8pbO5HXDi6kkawaXL/csCT8mgmI5UJaFU61pD2Fg6o/Pwdto3/f2YuDjyX
qpOzITwwuT6QqmCoF8F8KaRNjdVS3bB62VEaJYdtz9JL3KuBDapb+6wFdsUmjrv0SPbqB73Woa0w
2LW8ZqCbNj9CdzVnCa66UcQBIe4rfLLwEciq3cz3WBvdxtMrMHOd6rvU79InAR/7sntFb4zVum5g
gjayrzlNnz+gzVQknL2PRDAJqEz1TqXCLP/+x59HmcWgLDZ1FHUZ58kRZkAVLVXLI+nfqyU2rlJ/
7RxL5EOIvw+mIUH0VkF6Jb2LvpX6mpkCFbtd4SJnxlL6Tk56GI9IXkO20lULKgpkCQWCVoH1uGIY
S0r8Q7vBonzHDxRuluLKbGZOdsstAfTIOgZtn1QsUAy2HZxoz8i4RfcnGBV3ZdTa/WKOGJynEzGq
bVVnalu5rOix5wDZ7Kgsdc4Q4yKnYY2LdXxg61KxOHrgCLqWr/8sdlOOKJaBhQRxJgEEs7oQmCG5
xyvZAqnDofVDokLK1IKUpnyFQFJUon6lj3taRULDxSgnL3zQifmLVq+ysWi2IRdgPGwxiaVnhbhN
W18SddmztD70nQc65loKHIncsCj/bBVUG7xRF/jpwyw7kRzJvi7hrxB/bPObimh+i+dxlkrrV4Cc
MdE+4rC8HlIdHs5CPUJxom86DYwBnTxpGVr5dvBzdnfMjAgpAFxQGZ39jiDXeLRP64Z3tkvNyCVJ
Ns7pz3x354qLY1mqN12P769jYLW6aOZp88PC7+p0KZfBcCpoEC9WSfTajb80mJy1TR7oEUJsQ656
kUkXTeMPelVLF/ENcG0bhSKNulcplXFHlAZDGolTpoBZae4/MoSmAwwjL0IxOV3YCygn4Aj5HxnD
Ij5prsvg5f8Ern3QOWQpmW5Xlq6MY7yvvMpA3v9UWTzfooUkg23H13+hOGOci43FitYDS79meqMe
1PJLmGyOnJTAlTzzQv5oHEDdpWUUdmcm3tnauPMPFGAhGncb0zF9nexsHZVgmVizilvk+tw7xSuu
eBJ7Zl96TqdEyqbNU2whJQIzEVsZL8VAvNszSXUUT59cN+fetLmZUvHusQ0+8dkksZOOWPpCL00T
qxyqVoHmlC8YDuJJg2xeEwgURG5S3SZlEWoqcUe57o6IwApkN2wqXX4k7L8Q/d0sKDjAXKClbs2m
WffsSRRc1cxjw8A2sPKhSsEQwYk/XYktqtC3QpP5yu7EjSqLd55PVaCfXClKiwqO8PWoswFpzfT7
oH3mFhklixueScYtOnhB2LvyBJPzQwnyHnJXtTGdX5VzDnxHdJKoMBowAf/x1OkwBR2hhBYXlOTh
tgUOrsxzVjKXovbSQBzU3qganlWHyHBrIscYoCjgXmJOneziXF54CK5NwNG6RalyAsBXK3hbxmsq
CTMMx45mnIZ+u+uTFP5Oc8+b7DILwSNOkMt0WRi6NDrJazNpwFUzwWNmMzKBdfexTteA6FiJ49gh
cBu9f7xGtJRs5aOi98DD3v0zjR5TLM0waei3/hMXhmdQ/g8FYyhG4zjNGM9FNm58MiqJPlbVt5E/
0iT42vO7CbVBN5OgSE3m12DGcGlUIIwLBI53jF0oXVivyQHsmGm5erKjNqEXkRFwIM2SBVvh9013
squy5VvRLYFbt1beXYvdEk3SQmkyCFdFeJGiTaLLbYNJzgfQWRdlmCiBYbqKgHIc03WQ1oiiJWMq
8MQsT+mFa8g1LIL2uNPUiozyKv+ZeXO3QHxbWAHVpTOzECSOKo1Blj0WSZRueJVxKXRXHR4Yh8ex
90nZyqwb7EYfMnvTGRGF7/G65i2kNy9JP8et7JwGZa/oSqzeYvmsteu1C15hyFU5NUQoFE+o38Vq
y45DeF8rsNV9Pyir0TZO35b1/KY6d0guWx6YcgoieHREsj6LhHYmX8ilR8BrkNvL7ALM+v0258T6
XAnibhzkDCmS65HkdlwAWoihanii/KgnajBx/e4MMGpeShAHCaxKZncAYc+xilNcvG/KjpyJrJM4
z6lnAuAh+NXNwtBot1lL/NEvy+88yt4gmTSBxIv4zig9Fk7ICtHfWYZrIkUYqi9eFzYdjg2JoHOk
FLJPh7n0z8V1Z8V8vYBayHwOitUwfPPfnL9xQMRvLBUf8lQR+bpI0ZUUBFKf+cMcHJbrT7YyOeCN
l5eacOF8oDO9xJT7YAD6HZ34IY+P6q9c+p2fdzB9GWyc9S21uJ25X7Brml+pigXhRU2Getj8ftl5
z02INgoMANQWnrIY1GM4SA3olmGkphUOkhrkDq4QtxZ5UyeokxKy/BxbxjW6TcpW78rzcfFGQwZ0
eWHrM8pv4zW/7gp5U8qFvkEVKRbBYdScCqDU0JDGo0WNsrQ8W4YUeiN3GDjwI7cqFz+QPDWlMclp
NFgse/wP04cyDtOoyObJayrWxGQFtNzAyQVaEY7eixQN+w+5EQYqervAEvrgyO3xDzmkeKdPosJn
C4T00mpPhqkDBGIwFKfyl2pKFS9QqjiowMbUH8aG2k0a5NQ1TErX+8kJQ11ZgvVaBBoOyJHxvikd
42lLh3p6lgnL/agmqzw8Kc/BFpu8p4gbF6hNfbiUi0qIucDES/nAEtDcADiceHYmI7o3xYK4b2e+
NuymjbziY1/GjIbMg3nYPDm4DlOSmgsTxo1jAN7gObeMfXiJvboPb8EaqeiI0iAciRTqwxoSVfaR
jKdjZ4/C5UJS7OjR0O/i0gT8WLy0WqCUlWdZ6RfOah5i+11GDLcxl4gRsFuAVi2OBETzL+arJ+qU
f5R9OSxI7iGoSKGwuSvp69SRJOOwHyi16NPiltylgfC3M+8RMEP9EzIi8MBxT76xCoRiYSIhNXB8
oaR+fP5A+Q7XoINokqLVJI8WN1al0+qWxNbgOZ2sfjCeIJPm8LgCa4BTlE9mC2Ez/V/RyBuy7AWG
A6w7JAR/KOHlHbRnLykX804ApakP+oeUCkdgqg7JqjNjLOslxtYovbh1Vu2C02bLMYpLB6gqPRkj
CYmTFEh4yoWPdz1XFpoL0yktt8L65ct97gs3bQJnoLrVTs47CGMwyIsu5V9qDV7msxBq09y1VUH9
sqTjKuQM6nqrO7oc82LOlUr7LmkEh66YCkbSpZjfWN7jtKICZVc2HXGevdbx4bQPVioX+JhFJ0uD
yOpaLpNJqtjKSk6JCS/EJu90fznLKlzb16d61ez+08z1iL3y8J/RKdDbG3/wakUmNfwlKYjgc6Y3
Ckcjcgk4k1p7GR7xiFrk8ZS8zLLaTcnRyMa2xsD5/qrjeVOUAiJditnRvTayBXBvYysD4hBZo8HK
rkFGJTFRuAZgvbZQTtgTCqKyMTLmWHg2z/FmAFCtY55Y2mWsJLMF9spQs/xprWS++w62hG+jWLPn
JpdXdGWGytUMMXTQTM1JMEDYKUwRO3nhUBMWiWcimcyAa6CUf4nmB3EcWwCCD0qMsqraw1E6q4d7
7oDlrdOtTKY7rfJ54vRp8gkMNZA9WxtFqp0x8enTPh+D4SkOu1cLSJoka1uTDLsGoGG/iIrMzmeQ
VVtyRW3MJL47KPenMQAGAXupXuAqzeOoTAoxL19toLJRVoWAeO+Z1tKT6l9aKdYqSNLB+u8FqMSR
8+VadRUpALEc4H73H99CdWodAvPnvs6vvT1dNPhWE1x75QqGLyz0ACHV+L9XP8ICiCZxUD1uR5DI
y1/mxfepiPcIXTE0cG6G21I2mNIn7dxyZujMw9Zmk2BpND1YLTQhBwnbFijWox2LLRScTiQgKKW0
j0XjLK7PZyp4QA5RMxBuhvXbMgyAgYBO6EuCZoXigBNAVQ48Tu8csIEqQ2kmSLG8EZ+VqCXh3Aai
1DMry90YqRtNxe67KGDPr2NnVTzGSu/+1len5DMM+dQzVPIA8qFk36h0ApBnFSeVRvgs9rIPqGvr
k4pv9FI+2ylHLIyHnQauQpIb+MO+6pGgOvfzehtAm49K8vfe7KzFCAln/GqNH1UPSepZAEWT7soX
EF7tV7VxdqU3BBTa8K+RjxmSmlkE1uAzabz8XOpf0UUDGSprV/GaDJijtvFRNeNEwFqMR9IcUvvf
Aj2wZp7N7UOsjR69Sb2c6bXW7k6zItwZyyh7vX2BmTYxhBHAzaHEN7p+BPZZmOPAe4ID/QIBJRKH
Nl+mTzNnLaJKH3FA73obRK4Tr7HYSFOsnU4R1QpXy2IZgwBeKjMs7GdLqxRkG95/9LWShW0C1jIh
PFAWXjFsfZJAKCwrPnqjwEodCW+DGl9X7txh+f+PXE7lQQpQs1VMSsjvFctEMArk5VPBQ10dSZJS
6cmjfEDYGc4tlVGxEbsgJ1ZBYldFA5Le21G1avbH60ZQ42w/WJbfIyDwSMdKbHtNhxIZkegFbb1s
lJAEhL/05n/Qv0w29JRfv/NWz6KY5Lo4ip8S8xanQKRWOXGjDnzcQA5i/5k8t7zz7KENXx9Sb3wI
Jsbf2/o8X42jiVCHCZNdCis8Li6pl9FWOJbspIPYVypd16AHqcbKcc2Rv5Iclu9XeC0OcHRMJ8DP
+t36VLa1XjX807qvPoV65EU2DTdRnzBD7BL+EYIqj4Re2EQ+EG+XB9hUiMrkL2frZX4Jr5sRAZFM
JF7LyIuNm9UqLCRZyE6TbtSzd/9BUsUrNjICMKkQUN/AFeW6moCBOs1xLx6eHl6lbIGZK789Ugfa
4b0Wg/VdUhFl10T4P9x2qCwK8AvMc0GFg8+jWKLnwyyM3BfhcYcapfn6lhAPQCnFwi+oWBjlnULN
gghzWCV7XgtuXPMsl0YF28KxsJIQnRn50TneNZrer1kli5PvgLDll1lwA1iKc8ErZglIzLybARbW
wE2MJAwwVnAfJ2E4i2VsrO1pZYpF4bGvQLXmAFFixGHurVNicoxM8hUZJSdc1NYiFiQWRpMh0e3S
gJoji5+1IN15W1y4IePSFERtTDxeLrPOt7SK7qeVSmBorzdr/byZYY8+LAas6IaiDJ/ICNkhqu1d
wuLebrIr1k2CmqZOHW/aFoz7/W5LW/NJ1cLfLPdWAAPE8f1AD7xht23N5g5AZ4fY11FjIqJflbr6
B9Kr8TotEpVJnRqjYzjgDDCMFJQQyOdmoxWpLcpqe4OXUwALUH3yhcLI8VT+ShoyGZYSoE2s9a8L
n53jLYR1n5w16ifFmhx7lOBM6IDl24gH5nvEHmxIYbMyUxIANb2iFr1tFxQ1d7HbQJWmgoAE1BeF
NQoxU1d6DJoSwadSdIAQExfjn2cgKpRZ8trNrfOkl3Hh4pH3xMDwyWyRQCH7Jz9igYoKfYXpmmIb
vSEVCcANjy7PJ9a1LoCbrIpjaP96kPV20Cr6X2KAXYkqJPX9i9jn092A7XDXeG4w2vxka1PbsIbf
zN1KlC/LANrdZs0sy0XGl2fBWIBMyhlAjA2YG9Izg6b4F3xdI02xuWqy4j73dfzZI2reWIp7XZ/G
9jSxU0Q+WIXj72r7aZY7C4zDFhDWYi67En9BixPIt3HYOw8Jt6jcHPzCEXdMD1g+NT9N80M+8GEh
6Z+3I4HBdbxYF1upb5vIxnmaQLOs8GSxVLSNn03ehlRtFIScY0BgLyycDF/T+xy8DSQO6tSsOpPd
yDnHoJwWpnTKo3nDSbOiwMBkBLZ1mdPw0Nnhf6J/Xe/GGpBXO7kMPauLhBXB6suLOVVoALZqGsKR
LhKVEtP6bVlCXArw+0aad+FDjAJDJAdhn3h12DSCI9GnJ2cdtIznmUYVbPfPdI2QwzCgjCDEMkRC
4v3ccHZN3PXKN5wo0kfumtLu7ZWPlGnKiJTb1HSmJ4LCokBRjUzO+T2mP2b47HTMqP4rLJ24xRUi
Pwe8sDBCZ+9zxqDOAcBrAwjL4DuFKNSoMlvsO7+jORKhPJhLsD26MOMMRMp2fvoNJon51bpaIP2i
6HD/ascSTf1Mqu85b+FkVMeqxf3B/vWAninjPyqZ7G9TAmBKS+Gmf4Nsul2TShOa5VHO2JkwVP46
FOTzF+8+zjT6RlZo0SfaieBm5byBPoGdtps4ylnJQ/+QJw6UmU1GX7YltdLHgYsMatNM2xtvKyft
kgj5Z5dJ3VTpNccwJFT7OmX3c4ouR116bMeR6r37MJ6+lAC8o+mCcRM3ZfLURo6fqlOdWMLjDp97
h07WmyNHeDoUf6OZMRDf80SnmYbsgQNmZNg2AXjahBghbp3pdDwtlj7PlqBSrAJKACMr5yOmt3Vg
NDZNOB0MhFvudN+BX5h87CnrTirymipkDEYhji2AzpFtlWlN0UVIC5iI84Bkt6iIJ+eTMNIj493X
TNO4OQ7E5J8O2r4iTOKm1iSst2cyifGnIFnfukw8lwChWrdUNH+K302kdpPL4Y+0PeiNV/uwyDIJ
DOU5hDJAnvbsVTDNuTpy7r/siSneO/Z2qoQPudi6UjSbuea/VDl5eYB2waxVQjHHtC/hAGbvBjax
kRP1iGxGwryIYKOQ5qqAgavlNZlCcYKCHOJDegn5Neq6C5meC2AWVFsap6QMRcH7pP2fDa+GBq0a
3oHbWkgofGnSFYHv30568GwCN/oSg7cVs6ulUir/z+wE3Ef7Ft4bTS+9DkMW+dS+67f+i4yPTDwH
qPXwA3H7hG2RpP75OAuiMSmvMTD5NHRjwbXOtBmtht65PBZspgV22eFm9yKTMLAKpWsdfhukzztJ
DV9+Ppas3Qq/slYmAs2INhm3Ix3TuFpJoFGhfpkmFK6aQpk9EB2M8+q5A3SdxlHvxoi1+1LyY38a
H8VfJngriHZU+MsAAknuMx3eX7YBv0QRwzib+CKvU2H1TuP22G1/O7b0P62zl9IJU9yaXo3040tm
LvK9eFSU/zQ1IN03R4jAKdr5yULlcNvKLjSI+5/mrVWYZ4RphzcRWndbe9GP3g+1+PumGbDa3I14
gbg+feiUTKAZRX9IRuufGrEOLN365at2noYyqM0ozMTIe3AsoJ/IkJC6ItlGKZ/HllPw6aeVdyw7
b+8xOiJ9lbZg+pHivCJ4ENPalvITlEsf8FKg0+D9Wt4IGmRfJlPU0d6+zEOoPgBJW8pYjksFrO5H
G9UIeL01vVWTYJIZaSqq27RoeWFaDJ9FFFJ6BI7IbragC6IDR84KSL7nClT/Wc2sARyehCfsOSEU
gwlEps3Exrn7aAVqTmS/yv8o5r9nU7s9yCqbg05y3gCuD3NlNw0otqbGjo/g/3JEThCzSZBZ5bHu
HLGTLSteAcgXwToMOGdn/Q5H+8dotNh2IDhLbeKzd87BTFXJmy7QXu/bT7jKq3tq3320MqSJ2k+5
h2h+vPhLwsWv3cWvEjQf4qe+fnL9vRMiIzmkvIACJbiROUx8xHVck1AH2EA22OaKstxi7LtpBpye
69tltp+bct9hOGMS4aqrs0RbEy9+KLPnf2sgAAsHsyj0LbQnV99LVcY5qVaVHrqz1OJsAKa7Em/8
FdZfxRDwqvsqba4b4W5y3QDS5qDiBwEWJNKiOC55TscUylplh4KZk51/U/vUtzzvFlsnbU0rpbv4
QSWoJ83NM5sF++1vqO8r65N73lG02uMPtRIPv3kXidiQ69NTBDXgS/93b7aXqDWPTWbep7vwYvB2
hmgEs20j1LxYAPfF7AjSxT2xg25XpmNxMXVXruCN+lOOpfUCZ9NemRFWguciSTNNDLEnq0DhLCpF
yyZmlixD1o7YGMPUzhRSSTLVfLZQvnVcJrU6T9Rwc1uH7gNsHg4M31D/DqKS+53wEpHhMiECBzW9
12aCiUuGtANaXfE6KgcajjXzSmQuMtACMxY/V4phzKNs+5zAlLtLvzTFOdu+DkNMSdMg5FOl0x7k
IFa0x0Bwx5UXvDk4S9uc7OW+QTWwSW9R4no1b3//HHggq8DjjzIstVN4gj7sWF3hcyhZSHC3mF0o
z/mKuByZNfZSxzWHqD03N8Lk3+Rj4hxrSvI0Yi+/37ltcT+YVb56YihC6CCaioPVpKDBBTod2BZa
m7Qg1E7A2lW4qygl5Mm89oIU5r9ytUuSz5Jtw/FzyLhrHZeTULZD8jW1VHmvoPGFrXSBV0xEUMXh
6v8712jiimEsxkn5i398uOUYpIjdvdRELdHOICkhBlt7D30DoXWL6WWZzCG3kC06FYEmMdCUew+X
N/c7KMPy7C4fEWEwvKrxH1460S3m1Wq0+wt26cKosmPHxWgtGhyUVZelYuSl5wwuY8eZEtnjyy+k
qkjV2/C8l4MlX+uyN96dl9M0ntxsE05pokvvDbBjKEb1LwvqbZDEe+gnABXiXcPYBsSCVoC7j5G6
YjtCGDZODtBylYQfjgnx/C1FRhH6wMvLrTIayxa/PPxng3N0tWehOsflAHhPgyeKt1hXKnZtDT7E
u3CrrhsDlWUnDQtkqYHtVcqusF7rdGtZZcbe+1D3OGrBB0sGWMU1R1Jk/HI18mEnfvr0hZv0NfFC
Dxo2WqISVgdQyVuZ7jPBhXXJV4ghQy17uPCXGSsWhSJpZF8epV3U4MJxd0Wd5ggB91i2rwpDo9yy
0DLlzaYUeDD27U4iH5GHWx2teuOxYEFjJmucTXK7YwFPywpKc8Imk3PtdKsHRA8pj36hzGhpo0xx
nlVFqo6f7Zrqew8cACPLNWfnTBiDh3QGDUK4Lr+2eRczJ0YiTRtmgBQHWfr5KeFXjOCILZVBxACS
4NiH4a2W7mPLNa1TGpoSl59rjegkMlKsDgCMr4BmT09RvMOvo5414ZdTJl2F17sE7zcg5tk+SgXQ
cNKhUBdqaCP9J/iJBuCnwqarIb+FY+S/tTv08GU1DbJhHTlBGcihLf7M2D3HL/IF4QxIpzHF6grv
MDAuY5AAxpQFp8fsdSLz8K7XsQ9BHio16DgP8lAIMvinhVGgTzIlsfoGx2/Tq650qtHhDhxEBLzF
wgcTjC0Ye6qCWcRLYx5hUAx2kjXxEiipGQbX0E1yQh0Tzb5Xh80PA/z2/u92Qz/x6hBFFubD6+NP
RnzTFgOeZEaT8hTM8ZhFWO730xxPEI4lLgfe0OkzVTxYa+WSTiqH+J1DuKDxcN2Evn2qAXqXQwd3
0yoOHu7xNpmzCxRxF2I3d7dkslJf08DQ5vLbxxqEOtBGmF1RaFsEOzVOViJHhzTMtPrWgHoBWbNS
9QDtYQIogJqmJFZAx47Xb9V3af0sU7PxKYMj1WFfhJEqoSvwb9Cs6EB0nny2kMYr72BDqSZ1P7j0
C9meGP7CNMohTWMMlimWKRfpNkb25nbSuRxf4HsxtxV9CbR/s7Ix9mFx775k0dbHxDVJKVXMdNvD
nPq+WxBaf+2seqOTaZIDKwdS/v6MjEH9R84Z8JCi1kY4qIeOnRm5QYdp9ZuhPz+gRt3IOWWRisnr
MrFy3SWAlhlD4lMDdsNrzzHjHfRmb1QJkD/J+8rub4grr3puKcI9YbyKb8J5Jr3lPjJeoIGE6pgo
M+09WdsuLwX+5ZYxBUeuUQU3ImlEIDWb+mxcou534VssD8EKyuzTynuweZemptx0K5JPX7yuB39j
ejfvxzEr77j9EltrcidsVmzJkZ3og5MUw2GIXHkymztNt9T+XflSIxq1PYEsN5sxx3zb6MWQ5pch
3dqyo81qIUWGdk7mmPYo5VOSX/Z7qQzgRa54ItMPE/93JxHmdrmklfwkV3dVj2aWLYm19KWG08Vx
V6kR8xkC4LPCt2YvY71N6R8BfpqDZ/bStAkBUNbPtn2tXuMaJYeeaCKlWslg7Co16UnDgasS6n+8
VIQLLqIwgBYsdO5CgCV70rt7WgcxUdLMWubSWyC7W6VbxYlsnL1lr6mURLsOcg3MPHgCUGk+yGbW
R9XamOrmAsl+Jf0/XBdrDXzYJzAJKNJMNbIeE811msa/tFsFiTrxt880jctj6royq7OaOFgAZ3/X
IW0Qz2/7mi3nclfUOnx8pdGq+PXlRxfSQP3P53hYmrdpnhX7Sv6SU0ph+LQye8Q905nfpJOpt6b7
jBI/Id8xjYJw5fhMKOIdu1DEi9qVDroW3armRg3KdLe4Mj43nW0e8y/PJV0TyK2a4A/ozwTWXTkK
ylvNyXnls/UcaYL0PCU/Vkef0KvUw68wbOykSXhKPGBB1gS/nWfboHKTYJ9XRWFPAVxkSiap7mqN
WKpYHLkxoitrdk0BjSMOO+TUj8rLMzYgKQISe0gNRsGI9NIGe7tLIHiq2rNxZ1A9oE+vGClFjX6o
aFKUcvUb/u3ICoqMxirDDhRH1iPu/J5xnJh0EfZd0mMaff3JoLETbPEzsWoiiZSTV57GmXkkWWeQ
vDLQRFGoMIDb20n9z0Bv+Sjz9CG4P0x9SsVkEmw6kBKKqYsFPDnMc4czJJWy8hW3giwC9yj4gCXj
nXMEkUu29vErsegLkVTq5XLtNgERbd21lOBOldVjFyJa+tQeS9N5T5cE1yyNn8sHrP7PGeqKrQ60
sLpg3Y08s/ZsbFyjmcKNmFC6n++kdXKxJ/Rp6hFNkKc9issSlVEU5w3mjkzwgYwKtGxqwlqVZ9xe
EjvUgVqsVfJrNKm6Af9Gz4xKyeGh9slA8Ou7pE9tBH6g8uHBu5x1X9UVcwNhccbl+JqTZDKcIWZ/
Q70LgSAxa7XFTjW/rR+qkncWGeNDsjs5bcCHM+rT8Tom8Xd51hzI8/1s5iL4rxSSmql8uGrNCx27
lCPHdVLx6VLdHTZvikQmqp5TJx7/Sq+uWuOdAMwqNJkQDusjbMeWDET+H3QN7ViT1/pccVkW5rhr
HIzF62HBM0+77+NECEpbVh6ytpK1CO+itjvvge+30tSAJ3F7YHYPUjXV2pGtiSbphzWCacF9ZIr7
XfSBoZakA0eKHlNOEffo7ijR4N84pf/d5bQNNp3LHQ/dAuK+h8BaQ/HASnRu81If/97HoDfHyANI
ZRty1BroUGpv9H6Y5/MKb19M5uDlX5wd41C7VxeOoMu2vVh6aIpDrxA1ujSTZ5EZrjb06KgWPy8s
AvGN90v6kXpPgGFp9iEIzgQQzmmwOhiZCdZZgxR3r1d6NbYguVpxSsb+KO7qeQTLxgu2akNCfOb1
jaDNPJU6r2gKmkPoi9oIiLid1Fa1liz9tgeyQbTsVINRrfnqgZT584xl4WWz2aIgZ8B8fPkxRZnx
OfrXPkmKd/aZdRLyKp7+T9y6RW+kz2rDdgyxWdWSDkB3+kogha2ainkHK92EVbi3pgYOTlwcoRTy
zyTM5ZJmjoPglvI19XPQKqQhnKf2usH9Ne5QIaFUCsbB9SwY8J/LoH6Hd4YofwH9zHyTSTLn1fMX
vhOMEKoetAqwMlCP3yOo2uXP33PKzzD56OLVoQzd19kFAERr8o1+PGchrY9Suk+kI5OBUhPOOvuk
le9dxbS1z2MQh+YCqHt15JAr97hulDEIVIyeHpkATZRNGoO6yGmjt4dQONReK7aoMLxxpoAnM4+0
vprnjiHUsazMZtZF+lU4XP69EukT+qgknkNBSGUYOflOUoFulicUUwfZJiy5gBWCQ/jUjiujNmjT
QEjok/s6pXM4ePbn90TGHl/hfoIlyKpMS+Z/yhCJXIDIoChOVIbWbfwpdeQbu1DwshhlZppnxL8h
4d26C8HxuyJgXKa2PqVwhhfsBSHb/my43qNHbNQz2TdddV1Yuz6E03jDhbMWX+cLps9UfMGySVxA
y71ULozvy8Y53fhCR2mFjSU57b8pi3b1RK08Qr4Ix6NSteGI8kyey3Y0gxYDkMwPkwD2sjPZ/9jR
gtuC1NlrJZBnWHkkDJIKFZjxrZ2d58qPJmZKF5AE3P85jYd2xeHeGRo0f951oxvB9ns+kM0tRFmK
58KHquWG9cn3NXaud0HyeNJJ3B6M2uOKhI6cxtxxBX59f59thsjjcLpBbFneeaMM9c05lGvv1NEv
kykk/ojNwxKJ2uQJ9FpqHBnkOQtcm52jTaR/SnO5CPwSRxkPr81O1EHKJupuWB3khmWp1zsZ5tYA
8B1ggWpI5wxbBu57GAPLZYRMI8PqsWzuN+yxmtcB200jszWWmL1F915roL3JhYMxAjNpZ2RyWxaU
RTzMQV29Z9kDw1auKqwhSfK81PUtwWV2/LLaVTDeREt8phWwwB7Oog6oLB/OZt+Fuz2ZdPhB6aQW
8nd4Vavn5aB+LbbzMzgBbjE1P4Mye+kLGMqspM2DvC9Zz73Pi3YGVtwNnmH2lSchBaLfXeMq3HKI
CdQaELgwjXh9WycGyZneBuhQvI/jF/SHuZcBgZekTsK/UMO/7U8kKSyBrf1BhJgkxf72PuhzSbwC
/csvqKh3vOaPeK90OPZs8VdmhnIE7SJfiUJl7JOJP9PCwh2/g7hF9OLsoE6UBVEOtfShYPfWiEen
gfHQH/4JjcUvXaYayfnFj9/e18gxrEBrke8nAAfBwtfcRWfhIReWb+jCOnYO9h+Obluw7K4Lh0Qu
FSA1uXxPYuFnr6jGKkH5png+30vxKDq49g/jCRvkv5t+oj9yapMZQbs3cUn6agERgnLEJSUNhmCk
VozHcw5NDn5vHbcqB9vu+LdWN31gz0T3eIexBDjRKhffyvrj8PckkeojYWKEhttMRP6HF0FR7R78
mdWvYfuqi2Jhm8DYwH/2VM4K274hQe1J9PWvJQmmb0IyQK/I/Qmn/JutREOqhtyoZfZhS28E27tt
HuHesRuYsk4wRNXb0cRM7TYsr98L/KMtXsCSmzjTB4YT/xKoKsuzYKFNQiSuEOQnV+Mh4ps1z7iO
VxCxMhW5IjzpvASCsw7dECQsGxB556tEVrM/pS4zf7psRakMkYwhkr88y19LJSAXfpX01HwCUO0c
GrWLmcSQq75qCUToW69F/3jAOFHQ6/T4HY81NpNosIuWluHZbhTMr5Vt7m+4+GqeOqcmtE/JQxth
RPEvqEYJVnx4GtsUQ3Ou6Nr2ElqAqBI34Nh4PL4HWfYXw0S0kd05CmI6uRVGvMOZ8Ejfup/NrqPd
zXvFk91qkF/EItR+JUuyjvNN4bBNMe7CJXgm93JeYXr/DXce3Aj3SXToNdWRX9EoqaspA6+xu/gT
EEMXqE558dqDztZPbv65j+cdVUW6B4rgN7bWvDdTxa3odrcUCq4kD3qFFdRFBMk1dAopz+x/C2fv
2G4ML8lW6Wa5qQz/r7pZSDO7JhpGx00mZbEU1NObjqg9ewmea0KPqa2s5aDdA4KaPi/DELf+klaF
WW2BIJmpdsrRbtCq+1IOgSNxLC5dglbhhbr6SJftTj6bfkDOxAngr0Ld0kuQU97i8hz1/RsxE386
cIrWdwhKt3op7T7EB9gcY7RAs65fOnVKSMi7D1QnZ2wMY7w/coa5ip8OCst2ITOasTK5I2UAlEgw
qYal0L9y/6Msb/vNFD/VOrCsIUklg7u1ES+7zzQmurVa8fxXSNhH2y65YvnzlvKP8O7tHCOx1tBn
PhN5rDV0rF+BM5tFNpifxzymLXCnIKPPs9sbSQh5VtEoFrnBynTnNRaB+YR22qOpS5cxVzBM1Qh0
1h+cb1KYvy80bbsnoUFd1TOyxpe+JRmTi9wK62++5ddRItLkEZe2zUs/dxYaj6rbqEBO3uqdhL1Z
PTbFLtX927zHYN+sePkbK1jw87qzhY+Oweh536VdjZaIk9mo3jn3k2/gekE2sorPejFDhHZAiKxg
JmH85aDDtBuIBaQxS9I56XWR9/UTHQYNeTMUMjvJCfcnBLNw+rLiPCyufuChfAnT4+jexYAZUV30
MOQ8K88HjyU/fJc7kpZfeYrRVsqC8VYesxfqxYmu0OyqW6ZcEKxsQ3Fr7HiTkoks+KcG44X8mUiO
CeJ/5ipqm8c2fhjRVUEHY6ntHuD4BNYikHrp/OPnbXI25QkIId5/3XTxiSOIlMwk+kSXAYPFN5AH
fp6WrhJqcAKyujaoA+QdRZ3bLrwaoRKkADxueau7LFGrUjuZWjyOMIbGLmCvTgpLCFENo+nS4QnZ
S9B09m4qGqH9M7TXXvAsnRdklo+gGjhdwR+BGQcaAOJR21TTJHVE3UaS+1f0SVuJfNQYxFrlu5zN
FXNokPCMOolvy71ul4zXYHdYILQs2rHRovvQYYvhkTOTE9g2tIwEIW0us8cz7e6/4qr1UOgPHfA/
bHpnKfsx9VIbd7H9pQzvyFvFhT99PjAgHZSYM70u/+GEpGW5XvOZyOBdkL77/8Ihk3uH7PaVp0i2
7SGL7OOLsDxR3k29uuGk+qwxsq/iMpauFK6Kf1w4kdm90nm/CuLS8U5xHjB4HzYz3UxcJ6Hv/Eqs
1ywQYq6RGwgvwbN8FYV/RV3JSOf1/2Ga6/cCWH3JbjzkxrprzHcLLIK4pv6aTwItzzb5fXWQkgoK
KtwOCSplhUozKOlYGF8tYkX6wSNq7KaWez5aXLrWgAyWlFAa1HN8Ot8V7FqS8JHmcUZjtvoH1ZoZ
XU9lkpojLDzwwsxxHQ6Ul6nsw0i02dBCzWEfy7jgsJn3Cn9KO23tnsIxKFZCtfpW96UZLdB2DDRz
dCAZyFFFbhntqRYvZYquYTvrkMhAP+J1NYn6kL73f/mtHtg0DjZQiBPk04byrxSHzI2j632vt9yN
FNj1ujaNUdimFebbC02JrSzUUisAEVBz806i8lOM2Lj99jafW13RFoq6nNgponWwkkAqy3efNYST
jXiSE0nSBi5Qzo6n9XzSPyG7gDL/CiYvLNBameqeMNU55bn250jpZZVeuit4ssqc1W4btmqa///E
VkTFbh1JV5ggx2NW4Tvi/TZe6JWxNVE2FKvb/zEgoH7T8aAJy7T2dESjI7vIkR1eua8SKEwoUfP8
kHWtFHpLFVSarqXxWpdxsTFYr9xDs7s/Pvt7Gy4xykmF8tLstQRaSB/AjlOtbUhDxuMmzJ42c65U
HfeNxxEW7Zv60AGz9HrP/G82f7QGWoA+AmP5RPa/S38XEVkb9cNT96WAUzfQ2BTsiDH6y/DlMMMy
ITQcGFWYn3xJP/y+okhHrJhOABuFV2vPx2LUrOXQe/GMG0aZc8YOHFJIATUm9CdkuuB+GVtBdzDK
b7PWxuonVg3d/z1kKPXjaKYW5DzpbEAKWP8fudQBVwxcUOyoYlpu5/uI6Iu+0eC++3u83JJ/LQSe
e0cWuxTkFmXYobuyYyN3TXEXmj4glpVF9u6SHIWJWNAJq1IHckAVO/slODnQWyMXSKsdAeQLNkbt
wxWMnCqWDkNn1eBn3kZDyZT/KVdC01Rn6NimW9pFBXxHE0Xy3IrmCPxHWs6GE4d+de58KndwhhMH
/sqBRTBPG4NLt8mIjnTY/emjN1MqRY0JljDQXBFFzflRQUyyPwV4hIktNSABTl1Zg6tDf76cRt1t
T8Q7vqCSr1n3Hm7OUvb+KcX9yuoRwqxI9+Lwzi0sHaK6NH+otps/2H6wO2ipjGChkvYLw9YKokSl
IyzGnMFBHreN6XrDFoi10cRnYM3rlEYW+ZdX9Z8fJMm0xBRdwuboDHyRzu3ZFSKv6aO7nXae/Nj2
T1LPEGKRAZxPsQzp9KlMjgHkEey3plHj3VHaLrWwwrnEaPuTBUcgv1vPkCeHVpfWYHjDRjn1uMiW
a8z3iHSf7mcWQuwZA9zdwbD48AaNbPgUsXWO0cITZRGunzAEinqEfwwJhZ3TVVfzrgZLQFg2GhZe
ERCv90L8aYAIckQb/QU/YpEzXpMPrSjniFfkn7qSsLgxYSoPr6bC0ODxa5OMqDjnA53qYnF5QjRz
ZvonqJEBcGrAmlKZ5n5HSJr5ou3JARuUzBfPDQeNp1BXH2roJ7VC+wh5UNKjX5LnoCy03bP996A/
48L7a9G6O3z4uurK4kEft2GhEmdhmaCeLv/IBHOUO4THPBSZsD+1MAtxwuLKP7FB3y6LXTJlljbx
xp5CAT2ytfhMbx/ozYIytNm2gyoiQ6VuMgirxXzgePF29ewfnsEKlqDCcCL2GwPMNypaKsxad4mq
DHhW1R8k+v1Dm178lppaDeuv3lQWy9j6AraRGO5K1ZNaHU043Wl3EGwGfV1MGW/SYCgtCLmPLvao
phRCUQhAO2GWcDv5vHQPhMZZ2AI01PBHNSxD0a1UrLi4sDIMsWjWwRwLkiQKJyuQf+1Fb02e8LZn
7uGalWBSc8Y/DiA4nxtM++yi5NbXYoq/VUC7Ia+G57fUE/YM6+VseCwlbjvHZ7bOhEyq9ikqIYGj
iLETs/fmZNh+q8ze9P5T+4szil3S8mJaLMNEHmKOpYOBxdPcm8dalw+x55FIJEdcmZVos4zm1n++
sf78NEHkCumcPmfL8pIpt3BWjpu2MuS51081aPQfuIM1AelB+xs44ZbutCYkJs93G4QCzfaeFbcp
2qCqEZHEi2wPKfYYpfQ017a5tkRtubgihd2A/aK/FCK3+pHx1ZNZT6jqpXhsulhzXxvGmH1cdxcE
fptotZo5OU+z6LCaJNiFa9wypNXWW7UcKh95S0JgXcu62WqBuV3jSb6ucRLXsnNxP+ttu2qqey+F
7t0XjH+2X2rEUAVjjPhOaDVE1n93USfJVbkGzIE+SISjGiXJ4LLjPXXGo3HC+ToLLVXXiIIm/i3B
ibhBp9RITeM4/cuWBOs0rzHSuzwKOa8NhmrIIweLq9+R5nhwqZ9AwUvDIrwKT63RtS5yCNA9gk6b
v7MhqrlD0vE0uGTRplDiTloYoycPgy2OrQ0LqDsCiubcuDLaQDFlc9XjY4XsApv3qK9a6hFzpM+x
2F8s3EgSidK8H3jsqBgHpT/DN4g5epEUHm6xSr6Ai3NIo/A0adIRkdF2s/9LBRTQNj6Ka18yXoNP
jJCXXiOD6uRGbiRhnIBhTxVDkLNVVgXyINuyl9Tnak3/BGEtj4Zd/6u2918OKHvbuYDp50Xuq6GR
kKLlEkxfQzV1AZHTgInLUela42AC7mGAE1KAeyZJUBW/PNWi7HYn9sUloLssaFrUdmJeS5v3CfF5
4GSLPt6Js2RNNbmNPZ1W2ulzkryc3x9+0hLFb7iLsBFsugwSeeiHLnNhUdwUu29L4lsXadLRjg17
8i6kqnYrvHkvlcK3K5SxCAOILlUWDzbAmDEaSXobhKC8T8Rx2Z2K4WaXcDAYNZSx/wozr40omU/R
xEFUFuDpiYZMrKYCwnMHunEy0MKojn8I1tM5slLYQ2z2Loai0N4lUyH5IsYv9UfnXuZbjTh9NpvR
LAvcrZINrzFdqrGg5rL8DK7p/z87ndlxDe+WBFjdFq0ItPdvew7lmOaKyKP11F3oZWb5OQAdEK/Q
p2GsAUo+bOx4mY9apGpaDZVm6Fl8I1lWkBoUV7nSFJHVP8J6t2OAJDW7rUnvCsdXKQeCErblVXnA
cIUQQKovJ2iQIzFz8JFp5QWd63+a1FzyjNwcJTgnUgHsAvSys1r5SKqrrMiMcnWJuiU5MPNFhbhY
B3GlWb0qW+3MSoMeifPVnroRMZHqSYJBLGP0kcBan0Qmfa0WLkPYMfrZGn3hROXgk0GTIVSb8DZt
+RRH/FJF5bSN1c0uK1LKi5VUUpQIOLrgBTfKve435IA1hZEKBUi/i1eSL6Z9TRAs8XDT+de5l5T0
GxOxqyHbqIesW5LX7gtTAra7+Y8CFXlN7Bbo9LzzQNIjckkBe9v3SesBjkNGeOk6/lBvrfyhpgc+
s8GEuDCn5WL9xVDWKM67e0pw8RKXXJJ5Iof8AG7qLYW9Kb7F5488oSgB7tkULNDC5An4FyKQvMRD
XdAieC+1e00Hubw2f+qkdELXPHVFHs/nmn0NHuCqJdOSkVwuqYM+K2XcGZM8cHx5zMqtNSz5ms0F
GBKwG/Kl78kQlebVWfUAo2spGeTCuqddFVpSNAaLUe6M5LjZ+PdYwNCWSGSDXYrnV96h1Ax8bHBF
sRUROk49NBJIku27X/kinkYwAlOOwiLGLSbs5SHjP6a7cYEomY/cWVHMdBVY+GXsBNJf2kXv+l+r
DQnBhplz3bqpcdLhlTLhvMfPceqrsmIoWL/tJhOt/707XSFuuNmca8HXLqBGq4lTHc0tRs+Vl8R0
EQ4mIs8hSUBUv4MQZnlK13ZRSUfeD2EaaIWIt/qIrPTGqRK/Di0Vb8MO7SclLchIyJ0EKfCLTYnt
YaIOyII56ppoRQ0lke02ZDHRN2W7wjDGDXcrJORnCKGOyHt9Tu+yhllA4LQh2y2amairrRKfSiMu
wfcs1qBTx8M2/Rnrr5pORA+GQKcjDCke54KjiqCC9FC9YV+HTSBJexQAbAQ8zhKwbfI89im641Pq
mlpCp6O7zqDrwDQRMK9E03DoYghbaHNBU+Jl8n8anbvRUvjzaawWjFHmgXWmtpo9R3KvWUoFcpOT
aRLGDveT78uYgpyDCvKxSOm+z8plXFkG6+DImoxrN0n78XubDv7cFL5ToKenkGXuBGLulCGs9cFG
NszxVLhXMWro8yTHwJmsriMqtCIT/k4w1br0qhEg0jps/5LMRqGBHm4iWCG0PzB2A9ZPxiigobZH
3+gLUKOr+EoH/vaa5SMIElO3bTAekHXO9cewzPpoUDrIB9FKaiG2fg0UFduHMdLAREdlbRZSZS1Z
yNnOTWbbTDyRouo+qATLSHVXkltrmIKHcfXcsAB0J/lu4ZUZDYy1UCHcsIc7Xzg+JKjRDv4bszLw
Hc6CjEMXSOR5MLSpoy884c0kmKbPOjqFoIaU8Sp2hhvZ3LqgK0jRlD9QJPxtTBi2yjXkjwtjSB+s
JCNxIchRZHpwRYVtpmONLsBzj30kOAxuS6wrUvpRT3qhCEQvNHcFHA0A49ahdphTS4JWPQmmJxOw
XWlKFbIcjNrH7g45ZmF+9H2XOBF1K/9IUQcn9ZF6JwjOuBeY5nUuuqWnccs0SDnr/FukgeJrsQbo
JvBjxk2ZEBi8a5IqfPCUJeOj2JOKF/soryb8Fvnta6PfwZ1AJhDDCgxygwqoHmOhg7oCVWh33+Dt
5VU/C52dTp1FF0oMB0WOIQyj3ah160RNAe0hL6WcCgLLlGxBCr1W+uBOrY0PVcP9r1uaBYV9d8N2
95s34IbPWN1tJZWqAsg4fwSgZAobrkQf0e9KCVdrY0pbkUxLhXTWHeS/FhwG3mIcmBL1LXxSiicV
CGfvP6gFkmVQxSQQPSyxBTDjRntw1aDCb2Qv5+MB4UlTs6x5phW5VWkOkKF/t8E0NxRHs6SFGG84
BK0jSkQN3quSTHQ2/EN7x7Lz4STyeu1IW2vckc6D8EzSgn0QC7rCgEIvaHGH8v4W90awXl4icweZ
3vYZB4Z20ceViyEfAokM8vxs9StRxcBzLN55tHXTd0NN0L3zO34/2XZqV5xBxZUL8Fgn6ghyaWuK
Wwi68jxf8Q9NRi1hr2s+f0aMjXtGYuD/5Wgngdiyqk/Qz+Pywe/xODOJ1dZGogTvoKlWCX71O6pt
EaLu3RC6utDSnyKnLIdFn4QIVV5I314L3/eYfCkzCkPtJbgdaGGFI07nguSE6m6KcdCqypGhq6lJ
wHkNfGR+6exXhY5j/rdq+ZdPkMsPO/kLtRmZHlrg+MFlk2V+r+9qIMYQO8+hQvNxcWyJICAaJl5Q
c4tu03c0R5fiX95WZMEH9IIk0QfPbKOf0iE8xVqiE7FSDnkY5MmiwjQCTyAuA4w27vElhOCM0VeL
wcpSTlrCMNtdHvBXwnwSdwOPjZZEF6H8lj7MUvleBp1fmTs3Fi2LAc7JTSG/lcWh5bb0cY+Q9zqJ
bb8XzfL16NeHnOkG+r2dB4KHVl9nq4tyMAjRbSuHl2JoNJMH7rFAUI/014BCKv8ZxZ8FXoLu1OyX
1pIAKHfUvVM2nUnBeSkBWoGDfobLQyFNwNicwpk+UlEbWj1S+PQLGJjpzyBBUyzt/UPKBs6t3BkV
Oc3wi11jPqwdvOZekS8LSTkQs9ElXJZhFm68hopLbCaY1qYNFCaJi4C9TvbKq3Xza/1dCBQ9lOkF
x4lUuIQBLKsYe8rhVeeZowpYTCjZJiyjBrJ7TE3VSHK2JTQH6fYBKqlIp0pj6ZPHRFOGkKfeQPVB
FUB1utpnpuLCPhS7u4Vq0P9JxAP8OZWhTkQs7DU8BLPE6MeReyuqHszuma2cXFXmKamQAYWDZwQq
MI7Jj97i7hN1X+7TMYoIMnUuiuMISvsN4klhMY8oWK/qK6+WAVELWpfODnT/gjvPkIkUHdRoCca4
oA3ATmWZn0Sa+CAg5Pa9jLjKy6n4gzqzV4QV1+C97LUqV9JDS9GeatNghswlfHry5Zg87cUJtqpd
+sebPtp9sdiNol92BkKCAIE43ox+kDxzhonDNcYPuXCaJROMtB275Z6W6HFTG7OA7mrV68qa6FdQ
N9WgXvvtGsY3nOCA/30RKrXHUPp6hdRhqX/7NJ3OfoiAIcXhBppoGWVHWuUmnw6JB8dG+225atGE
FEf6Yu012u0VUTlKksymQYsg8r7Os/qmT9tAumk9HZpSGFPiuEV3JxsZIfR+krlJmOa7PCt33Jp5
RvIX9N7Nr4Xxsc3b4JAVyuMv7Hzg7u1/iTIXJQMV/6OZx9eEQXLCfAi4v2sUSSZwtIhoUJAnqCev
9/qjZnZjpeOP5l7CMOR8jXs/FKTStwNWCpPe/pnFZRcUgDnJFU2Fe+82cut0X4hnt0uwOPpw6XGQ
AOb+xhlxOfhB7FZCQKyMZRwB9FTTYHUDhIwB0VjKo7o+WX1uNMpOi4EA4go93Wee6bUt+HrhAoz2
KiYV9WdFFER2FdlEAdpCvHRDTBLkvYEGNeZnEGoYX7rtTTRvY35V1o0ViVpNAfDNI89EPkYkZtIu
sDpvRmb9IZ6hs5HdXxhMzL9QM1IenPouH5TRs/Nfu/wiV+wepFf32sW7K4CRuy4NP1pt1igSI3BZ
TP2oxXgWS19e7mpHHoFGKD/VBnBVVOyKVqty+ocHxuo2Mrbs0GPQ9ZlhLPfJMlxBCU6ZwQPFI4hf
yuLPqBS2/y+dmnl6B5LZe2rY7XOXnlCy+D6iHHXKPhJYNIpHh/QumRP0qtYGaGzYMBn0Ra2IjBPN
eyFQjzv/0KPsi99vK3dwdYecnaeqTmRwLSxf3LvhX7MGHrAbxYR3WXllu5UrdpNgKlSh1/6UnG9j
2silv3JyKT5TaKoZ+2L3JJPmGXxk71nmJ+5I2hCgu4mS/qR9RNW8GTIULl+jtnrkDfJEb4Drphoj
01XXe1xubvTcWaqoNfdE1Es8Ye0vjd9n1KlsmeFF3RwtrLVaw7zn+y6yEz/OzBlNvIgqvXhrsKbc
b2Q7H9tuvX4uM/LsWu3gOdMvJ2uHO6PV1A/Pldqv7NaNIcVz3F1oTfvdIs6J0frfRV3KCVpmhCo9
Sf61a9XtwuSVUb5yjjn4PwACE7SoQpllNm+VMAsE44B8dC8/HJndEug7qLlRrkvx+MdCU+Zhwhu1
ELiIh+v066Hi7mHBFPrRxu2wzWcdpjTERWyTe6TEO/GgVoUGCm8LzvYvzcqk9VDpXszdof5+MPqV
Be4t4UqUBkXFhA9iGNI0YOVbTIXuKZkGWgHewwv0jKrOnDwyB/XSCRL92nM8sY8QChkfnC/+ziRq
bHpGZieMHDBtsC9UH+GQe1bL+RfBsr1FQeh3EQDimfP3M+1FuorUu0/s4SQ+6jHW7QhEaa3k71NU
zrQM4yVLfaQe0PRaVOxhy2f6r35RcEDhKaOQcL4SMfGg7XLODtolU+GkSIAWdqm5NGJNa4qrMadn
LnMlmfUyH/WCbq1GsNzmpmeLtt/JcWrMR/N7ElnRzE2UVs+4103fz88JsoKWRUrtRIXVMGJaW6Sv
2r2YYhaj400W0kX6mjlej5jyC9cRimuf9LNGqfFUb3vGBIBX5i6r4lEMTL/T7yX5nAXqDRN1IKu2
Gi90L8aCMik1phmmHJW9TkxuVPAb/3//7fGkB8VpGxuDzfmcx99JTPdyFWRblRmoQdzSpWy6t5gS
rgX1YCZ+ZpMEGuIIx+VGqV8M0Z2kNohtQkU0waVTvvsJbzMNckX/zgceGE+LMBFswlBvaov1SnEw
M2qdpFxOCiZMprFco/okWFcJ/GFwPny1c/KnpR9Z3r5ksQuJZSfOvr9J5vISfQZyc1IZdLBckV99
FdXzNM5tKuhCzN/dBzIIoFs/61jaJB1nWWzX1ymyj30nxncSObOyudVLZY0smGkd8pJK2tdocm21
xAK0F7eMapBTGZjdBJCY0VA/hkHuyK5llqNVbeIVPzbrZa1+vVBhUATbEuHgtLU29VFTEPOe5871
Z0HA9YbbA7J46Tp1vOeMkng8ksJpzRphufEWNKpDedJFB2CkWLqiZPWplZth92QnqC5ulSF7qPvi
76KoCwOTT0Issxr8EE6BwBz43DRd2sz0hNLZb+syHVg6H4pITyvIcth8y7IdLFTetwMtWcp4Le65
f74zvKFbk8Hx/mIsCs5dXAo0Ubfr9+zbwcuOo30JEcTkFQt30Lm221rptWVHlccKX5hITU7Q8qpd
NPmMihCn7UQOTsBpthe5dXUdULoL+EnQiE9mi40ueCAkGFECXIX3JgsUT8MqHIhCidPUFzy7Ns5Q
Yj7Wt64O5HFOjYqsQk/PAjgtf8lPMnDJS/ufuwKXHJhZcp+XEkWDZs2Gnd+Equjm+0puAXKSIHTx
g8fGTE6BsO3l9GhvrZIQfctTRG2iLjW0e9oaBlbXtnqRBv1vxyiwYHIg4AQyYjgl7SZ3uwmqAJV3
m9KbPXJq6rKyPsaDUtRWjGiVKm0fZmCpUpuwUnExtHkvkqSKhs+lREUE+vc9zL4dbsbzZl1Zghwo
Ki+alrribUxZG7GZvKhlHDPmLzt0Xd59CCw0Zjt3dTaE2mlkLY+Z8eiOlhIKzPHkNBiFGdqBOIJP
ybYuHFgE/DLJ/3LALAAjELjecIsjgBETC2tOpcQxLsQY5pxXsMjii9/whvLdF38qWrZhnV7jQGm2
jvyiGvpLdQRHSaKEedePeFXeu1eL341EI+v4Q1YcMJJiFD8e5vWZXoQyykcOHmlKK7lrB9VqCxWn
c8f8pqpfTi2D9CvHv2h8ycFMR+wH4wF+g+thU4Ehc1cO0xm13yu60yfeRfsg26QPKRknQC3tO1xy
X5fGH+pCC6JSJL5DyhoBL6pE4zjQdYVaZWC0LCY/Vd13zs+qjk4vx/WaTTgF3X/NtLiH4aKBNBjh
H+wigD5ypREeuVJ+bkoYOZbOXxOaavjip/yBuDIBnBwttKTV9n5EKk9W07M66slSeUBn5ko4eY/4
8r320HWvj/uLbb8yax+ue5vGcgw0dWqsrR0JXM1c0ZgSlMXMe5HWGY1VsRlK4tCkG/7ytJ8Nd4Pf
3heE57/bK/3v1ukDzuVvD4B15A6hN6fUE5bx51xMCYNxwxii8R1q48ZVRcxOE7IjJKGVRft4F3JN
H8nl2ZoCY0zdp5qXK3lfUTuUPsgCOsBlf19I3A+ahIAB8sIZwIZYv98o4dVDvkeCZvZa9K2KTaM9
1UXtBC5hdyadTPomPzkJY681kVVJm5M5jZGs+OMtiWok4pS9vIG2nJ1uEnY9HiHelKkzSxn5XqMW
UQWgD8+hE4SBcp26A2JoEMW3GjffUYs7666xyDsxt0lggX7PzfLXnw90fatqmLH3XEJ/ouWx8Jbm
iXrkAQjnZYb1j9smijWplg8XMZrg4mWOYozos3sLn9HN1eWnQ1HCtcN7aFS4PFuUecuqIEiPSo//
034xkQfAR24gGgtI4A3/NQAfHys7KSEG0gpyL4SNeEGmIlUUz1+ZxDfFk6k+abTAd8oORfsJ1j5r
nSaL0x220v1WJCj2jzf/0amKYAojEZMPbJx43GXnCc7jrfSC9K3hsNX1D9nOzBR3D2RKx01QmabF
eMW5HiMIudHDKxSCnd+0ZM5RjPvRtl0InEmRukt0kHkSqJUMFp0GRomTPhqOKoOLgf6dDDgw54GS
jeZQ1vTQCLycIemumXv6PPxjop/yLpa5jMfx49gAaRGxSmCOQoy743wZPK0GpkFTuDfbIqGXKXeF
6ZkyZou+6Tm+FPmYN7IKwB55usbZbWSD5+j3K3e+3dqPIUKogr4GrmCWQ+MSwKAZn/fMhgKZ7Ecc
Yt4iKubBN+sTyr4t51w06Lr1QjWw1rhQXfLkqzFAOn99iuKSoZA+8sdf8OKrdU37d+ta/hYvdIfK
einoaCyW3oKsezO5bPA/b5VcFQMK42TJANUC77rJMXEaPOd8dCs1MzdYBorDIkhoqIox51sVRLUY
16CG6wux6kqO3dEcS+TLLkBEXKH/qix4BLME2k5wGXAP/kqf0Zfx8p8wLxOch4T5wtZSjK3WlHbF
qUGreIjlGbQhOqYVhEN41TUgLIcubUe1qHmih8JrmhLMuiCwsGQFlyEi4qo2UfFO9Nc7doEkc/HI
yzXZWhAiKgHz0cqY5yRTKEge4Se1xG3Tb3EhY6Dc8+bRJy9JmlpUs8AiKlxE/93UqGO0dBnrRT0j
uuRlZD16jJSS3q2QeWAPd+X/f5VUv03ks1sCyr0+ohiZpX4JCGTSkiCyhZPx2bI2bvYeXT/UH0bL
4t+9DJFQFDzvov0mhaBDzruIGnaZnyOtbMv6Jqr1ozbZHIlz6JmoGvnuhX2dx+l96+BxIoXiRUVP
DQ7lax7voMg0BkbPGH425iAoaND/bzPKNlsWJB/lNOQqi89p0Zk6RuUFIQH04iQo9T9xJ/D/KU4e
57uYYUg+0X9j8E+cNK3QHbKZ8uEjpX87L0zJLEFwN5aCBiGDN5r4PbSa2BWIz6Y+PW9e9lZ/dGpi
ORvqzQmLbU9c0KRZfXOM3CNHgOPm6QS1sWBcucr6Gn+lYAI5QLr1iDcW1XlPKujAuUyXX4EIlOqk
o4mhB6d3FC/XNgh2hut1eq3icR/4NGD1u52fKMs5II6RUfcplemZot/VCVwOQ2bx6VzQpsVpPRSJ
xtDNVAwfz58CRvlxuH0WAisKUboiGqd9uhciN0kMtW3EH90/nZKnpdbd+yM/IUM0QkwMTIk7f7nK
ec4t9vDFebhtDJ7PjmOSKwLSCXsnWiJ+9XfhepXuQ/dYPcMpCCWN99W4ritMXQQkeufXdeSL6mg6
7Z+/PqKeWGktC5VjwuPe3TvcKP/gU/ALI2Oye6YB8km2ddxWejOrfijEvxt+NxHfulljzsH0f2Pq
DcTCYDWgoMjPZXjXL3ryILvVgLRK8fSrWcHAe/4FonTrsmGuVI1Jnv1QWNRrKUw028JF7fta1LA7
E+qDot2mvWIu6XUgRO+Dcwk+zVapHIX7JYYBsFmWOm5AAUs60Sw8boXdVxQGR6PKcTItAhKV/08Y
zgL2how3ad3InEuxNSY/9HdgdWDijjc47mnV5yZ7ZXQadNLn7oRNoa8h/rDB+lPeu+gTUbimZ1IB
Iqx5BJ6OvAGJSECrlJPkhVAltvPENDud7L7ZBGFx+K8QZzK+8Xt5bZ8H/FeGQXGfdJ3uVu21sMAi
bEMbW1uqWv4UpHiMIDzr/oVZuMPi4yA6DdN0JqnVyeW8Y8rHV6UwGqgRwWNZ9Jt6NnTkh2gaoYML
sk0ema4hOa02neWZy+Z9GhWyvknacw7C6wsUPiVe0xz3S/iy/n/raOv8uYNoaOhTwKAkcwO7weve
1GqdiloSZfFUBVNAajTF7JCfzE8O92qhE6fYSTcVz1mCAUvpOAWdBQkfIG+YRDr+iVSBVLcsabKs
OCQcCYzweutLV75PJtBe6rWbl12NT65aYk2D0zGJkj8LfIEMVmLpVXc1qNvFDMT73vf0ssWWuXhh
PKCFsqJ3K9P+Hmkr4HUQVlvnEElZCDotW6U6K96ohTNRc4Oih32XHMTat+MY97tAjB9ybq+JVYCi
o2rSzoIJ1frhEATaMcfcHuGdfxQMJdK0X++sISyYKGeJwhzIv28UUNJADg10/hhRleHZJaoOi5Th
iAnunuFQQTAjwjSy8CSHlmGIu0HIr8ogufR4YKs5tSFQNjXfCzPooh3DJljfvpO/tYXNdrAJMzBz
vRNCDaPJla5GOP0cmDWdowJwhDpYp77T2CxiPMjVAGccsEIvQQzqUDb5ULYUYVc+ALmK32HP8JPK
3ESb/clgNVIP0RlSXXhlG75IOEzUzY5wbZeU1Fj+6/7MXYyQujsdZLNr2VqMtQsd0EXWxbDFyvHk
WP5rkttJ7zQPKWQ8gP0iGydAvEufd7Kaj4s2qsox+d0VDKBpBT//bkWfMac5tGbFZic2oHeXLnc0
wP6cWesxnezBG/DEk+0TY81hgxqsnrHa2mwBMwckPFFCARAo2gW6skrHNGKZMpjRhd0xkaANWD4K
ArJTtHLbKdxC1S80mDYBjWOXaR5JIWcSjkwFnL8DihxxDUo7h51vvJH7cAmPT92RBfbxvGiiRrzL
zMaMatsM1GWiYD97uX5/+JkkQ1rcj4SK/NX585iXGuSiclYG/ZtM/9ykz+GgZyUpgkcOx7HERWVu
KgXxFW0uo6y0qiltwg4YrUq+DYyL3ep7ofUwJwySZfqtS8NVVrSXDf2niabgwY/HCVKFji/Q432v
iOhja2uHA8/N1wBgDQXG5m1nufl5St1YLdPyS74mMvEl1uwuWyLBF7x7Dvxdm8lkH1AjsOw0nMXg
oqTVNpBWm0sXztjv2/qNCUQXOzwiC/JEPZ2+g+wvLef5Ps88YLT14ZNqqBQmlJ3QYEYOPmHSpW2T
9MBUCvM2II/2F7xopJDVXUYndjGem1Rc5pjdNet0TfQrPFAUDJ0AVTiy5EWm450+KKuDXUa60iWR
gCC3ZYoAONwXHMxRjPfL5JBhl2Yq7TbsAwNHEd6CbQJz+o1C7r7w7/hHXFVaOxV4p4uIkVM+W2Zd
iAsmtlK+tU9kFUv5CR8vyaMOslzLkNooUwn6xBGHe8IKLD3tcUHqoxgBn970r8lwrRGLUOKfcRUM
GstSUhGoZqgxpa8g1973aukhSNd9kBnwhmVL1il/KpbHcCywHT+WcxbWPsJwoq+4s8x4C9WqhfwV
egBL/hFs5KHdO1WVcbiF1qT8/5nd4ZsaJxqJqCz4Hf2JxjlM9BrRMCBegLLTi3OwSz1jk8YmrYiO
k72XsuwrIrwFnoN4H72L6Ye5jJ7eTS3u4gMUsUN9r/Tu5phCS2Y1olP2XXTGHSrJGn+rM3nybbO3
l60guU8WLvEpM7IHP1dXxebDly2vxfMoI6oNiB/yw2hG0h3tfcA2pzB9pzZukc+f1pg4KQ/WWCpK
ZNtweDJEkfvmJ/9AGeKz2tR3ldjp0Q1YOP3DhQ1fRAf/jAqN7h/fuB69NCMsOKwSkss7WYASEm8R
yvv68RAElphA7KLEH9vm61qLvndg/U+Qd2ACfazc8hMhKxZ5xX0pLHq8+Y/pwoV70hUB4KBYEsq4
SaXIIsAXbAFvhosV/48E2jIKp1BFa/doLAUcFK5T9zyC1jAOFFId5y0WHm4BiO3Da/V+R/zHGoma
bS7zWQ5b+DyEoNpxHifK5yhCgaZP5UOmYAuENwbQi+gnfkA4Ew0gKkHFjl4XZ93MlEvMZ6zr4gDt
NylpVEsM8446/1eFnzsc93xXEtPrHX2hGTliUhRArESghpE/gniTOO3KyjTKtLzrfR23nORAJ92v
LxZEJdDsG2UzhrGXBUz1+T0oJZVW0mNO+elfbx8DgsbN2gjMsBGJOYSeOXeOOBOkS01WcbaA+dkf
Shz/T+DLO97uLZDkKuGsscoepsYey84biEcC8V3b32MCMprkCUe2zB+AQjGJCwuSJfZcHwrz5/4j
7+NfiZSoZjTb1Knyxwhmyu1GIRO0O5lRppi8wPwumASXGNCFw/eROU5np8ifC9gg0J/K89Czrl8P
BGl70ejjhbZNSfpxFHWybS8HExBhVVrd6A0Cn+OF1EY/SsGnIXwgUINQ6O0PogmgndDuQYb1gJjK
7eZwSLZBPZev5H9HlRGcNclnX2S5DSG5zq4Le6sE8cYVzsBWHbpbJQFzXrwoei7EhRF7Jk7TR9BN
jizpwlycdYFTgGDIUHaPywm7zIrJrv9RnP6t7NobRLQ0SHjoGiqLjOP1mhuvjaukeVcOJvWbPVSA
jPuIL0bS23EsCipYKcS5pxmX6CDNLX7iRfGhhX05UEHPOE3oRyZzju3FrRr0NCmJtEehYCWrnImh
13ovA6i0/Y25y+GmHvdHR4lweKXnX/8Wvu6Y8J6aGlC7gTxD73cpM3f11yyxvuWne7NQT6bRtP4S
bJeYs89wkhjYXEwux/eIFp6yCf9lCRJfl8fJk7wwv0OB8YHJLDbg2KoC6SB1/9MRAt+YhCfD+kdH
7d7bdEAvrFFnNIiAbpLzMdz4+YvtX4BxQMnC1fP5yn64vy20azR2YfenVlemzIol8i3dwkWeIMPj
P8CzH1mxz2IoMRNyTFAYpu+MgmhKHGnK9bt1JtvzHrDUf1dJftRW7RknorE+cbLIJD8piDKF2Eb+
WQ+uBbQ/U58C301tYnnXNFqqmH6C4E7+w05RG5KztQB54NFObnVTlEXO0505bLtHW+8CCpY7er2R
dbEyYyntHxLPRHgEu4swrnfy5I2V7GFFtjaWAV8ehnEr7683N3Ijzw24Cmk19FN4WLQrJYwKobfv
G9Io9UO39d0HmomoUBfzcSVhqZRxl8zHNwcRAqhzVf0F+LKGE/kDqui+/Qx5uE/SrVuMWZ3kTTbr
dX7CwCYp2H6FuAR07s8STZL4ZytPNf9XmFzdIFXZKguIbVlBaCiVnR5GNGau/+vTGTDLhiCP6OEm
SToaEIwc5Goq/V7VGpk69jY2XFTUnOK2E6V2ghlku4sWAOQ7nFB/2BY5Rh04tXO+KIlFLgmeNwqG
hi2N077Zlkqq6ek6CWXMkzrygyA4TOJwVSSW03VL+ltg1C7G7j4B9wZUnLrcLb4jYsFHT4WCEEVI
bH5WT74LaBQuy0AGz+h2tWh0j/hn4sPt437tebHqWwjeK8OMuoQewQYHjKzUU3Tno677KARaGI51
7ByK0b7fQt2yYhgoxolZi2AOM45fzvQNy3MQVG3yybUgCRUswIWNy7Iw/AOM5jhOdQcdEnKjMgLm
VJJndHY/jvizZdoBjrb06Edv6TJjj59OpFrm6MvfTPA6sUVvqG3bT39aS6wLVwyLLJ2xzTTYsR9G
D6EnD5fipjuYV4WWfdviKZ63EHfFR0/YkCCXnARZQpVPzrJ0Msl0sPV23siV+qyseczlEQw4ocM6
ih9HiYfyvs8HP1HUC4DHfN2/B1PPNInI5G3J3keMaxPfHShNrX7v3et9QRWvCVMIGteekY+LgkOR
X8lEYXw0s/5ZXQhDDgzqE4xy6R1VOkOnHCbe3R5oldehFKX+2Fg7DNlSZ3XTIYL4VKsHkcULOi2h
hzYo8DKYLbCqCw4I+Je7hlkPrfEYbYfaYBSHRcWT3adqTua6fwso0OuYYpS1BdtSRipRrUkBIrS3
7bGlfsg3q4ueVJ0i2vRsBgRDxYODPOkD6O2IljC6nBxg1ujrwM1IW0sR24tl/x9CMQlGJS7MvAhR
TmM7DOOc/g7ZIt7sltjO3sl732zVfgzRD80nqmjV1va4UMipi4ftViYdl5mjq8X+lONwVTb8shFs
85xD/YXPBoLqHCN3NHsccoPI7dSQQtXexTmvUZT19aT+8msD4TcP/AHslhjvYbyLAejE61FifjiZ
J0sX9iSqx2hBFGPTHMVQ9VbOm8fkb2tQmoOsTyvCLpdhVnW8oNbW/3z6NiEpq13h/7wPI9DpRLqK
80DboN9izfaonZRTY28zIn3RrsfGih1kei84MzWIfZj8jvk4iTzmmHKaBivdmlHWKZWVaOdF/gx+
nL6IeAWkMnLWcDq1a2I7elrYoli/najPLLGu5z2/CwM2ipr87PXtPS0asxtT/7oh+1A5OCpLIXD5
JUhgvIuA2FdMAfMLyn05dRNHVC6zNUvUOZRelDA6adDYp8oioE5jduNJr/WrF1nR6d5cZcfSG/LZ
MwbCDRkzAabAOtzQvjwP/udKQs36fTxsbA7UncX7MUvVhQ3HSD/foLkZHI2EcqZDplORhLtnwKra
bBT38QSXkx9PL7uIC7u8FL99+2mjGAxjLBMt1qxBhpIM+p9koVaBW+zwiKmT7MJitFIFO72b7N6k
vjgR+dgy8WN+xfoEunxswkjtT+8twDckF/hIQSWE0WEoZzV8akeXhETehOtUOToz3ognfL4lq5od
yh2WQ7WBx/VYdzw3IXaTQFU0Z0/5jQWOk4dTHjdQ1tt28Nhdi4FZGcWNtx8x4uJTi5Yc+rmahNDh
hpnfnNdeq8gxaaCxRURG8CMJ9sUYKzszq7mUpOwDMmGZKktLT4fLOEZX4aPvxNkPuR1ebz/bf/di
XrQE7PnC1wNmXemiqqS9vwf/fX+2lPY9Vcktfq3J4MV07ujI8TEQ8RsmCfEHGheI+G14WEFLK6k4
cTowCRhnQ09y9q01xq38untIYArbn4b7ZH9+JP7HZ3scw8/csyWRrwAob/Ncxl9I6mkmG8fjcmeN
xmQaJ1/XjyYiunzFB9NEsV0/naCqAAI9q3GV6MUWDhHAGRRWJ5B3Yza2brBW3nXswpeiz+4Bd68W
tI1gfk9/ETnyMRVSEJfVjsXlJEESYeo2pWqcn/ryJFKbGvOy801QDuZ6YjqYpoFvxB0h03lNjUT+
r6QnXBmQyRJ02eH7GFXYq7oACJ4r/RpGr6DuTOvP0hdjkoq77eh+D2OQ94yopg140xPykmqnYZVJ
LfU7EVVaNDfd4ZEoVHPzJFS7Qdh0lbdb4hIorIm/5zCAB7WMoJmOmtIELf8i6/FXKJtydE75FK5X
fahF6O90hDB44R5ozBfOHK+/Y6lmmDau2EBSMx/uMCMw2vXGyKyb26chjvWAy4eMxkHm6Omaxt+n
+1tGSNiOIJ6p8YOalFr8RHNYhtOoH7qWcZKHdobTgJ8OlKlFxR3djLbkGYecD2M5QWm3s+akBE0a
8Fd3iE2Za69z0sCwuFZz7HPe66jeiTPAEZPeCqCvZ9DIiHtUT/qyHQ/uWq8uhUHNjXrP7E+2X5k+
hnrdlxWYWPM2eAQsSCObR2EhjXLFtCoW8Z0MTGyOMsCea5MdRcVM7tZJmBUQANwHVrmvgbBGOjq/
MLTPOLpcHDWEyszqrEdS6l9TmSus5oIKLZMcGMBWrlNQ6LTBRrt/AZeU1qTZZQZpJezOGktfaZ9W
PuhdqPH6zTrCFQon2b3Q7u5i0unwSEtQekxjIflDuyzvu4PdCCUjeDIkNlS2uyPjEDuWJssiO64G
2eIVZHei/roz5+l5KtVD66bwXpQJGuyAqmELJbDBIYpCcTLeHjBzI1iGehCx1jI/tkRkJCLfcObG
hibFCUQLWLjDmVMvDMVvhNNhozrmK46+7KKYxkdpDxDMy+MguTWMJv6rsGe7uT+FSY1UivL4a4JR
TUO3XGeVvzcfQLbZLIW/w0tQN0Yr0z3sbH4uUamkBtEX+ogz9xMfpt0mLwm4xcikITGngbrSagVZ
c0nP67V7zkqS+5Wjjf0s+qSB6wpj7v0JS1lKwlNANDTAipqtIpG1lDlr43LJ/rv7nBUtc3in/8Kn
3DLLVwowXKClMLrVmvoRzxCMaGH4tVh2rjDW2VchfPwL8xMh1bBOOHr7pJHpOxTW2n/DcjZGeSCV
y4TSoLFk+oJEPrcYSIJc0jPQ99+uX2lSIl2SQEqLHJ/XeIPmtGIA42DBRi0csuaztS61mp7rvGiz
U9NqWkMzuxeshJe6am/aRQvLfa3K1EB82lhGKadMkgIMvDMb91rcCSFQv4G48Heg1uvuXsq7iLS8
dcnSF+4TgeO88IMQa62PYIie6CPsvA/2XodrhqWOD/hzPl5orPjQ+ekx4JFVU4E5cu86nhDmrBT6
6mXwmSw23CXe34kLrXj/g7r3hQ2JlPS8jpH3/RaenqtH727B4sv0VNm/VOe6tE7jUiQ0rPInxb3s
USwfJE3CbMWDgxpapTVq0Es0Eh0pV/Qgk8sHz8trP3nE3MYPF8Dj6DQu4usx6jURg3NNcLdPnTut
/7GTpSzmkark1xkxXFd59a2t4+7uwyiWpfpGh3ceKdD7q++7vy+4aXiZJByDlMAQN1WI8f3YojKN
PddyDZ7c2mjdKg7znHqnBX0SOYnztbiWWjT9ZFE/Uwr5Ae0yTWTItYbWQMpSoGzmewyG+z46MCxQ
KdMTTbS+Gr8UUv/ZEZfjCAV4mcJ1CwxJhusxhzo33Ba2URRiAm7ZJWV1EqNAhyLQImW7DEW8rK4f
uT+MaFvlxGvTAUy7MyVjDDl0NGw0G9kl3R1Rb4dSLr5bHsXBBHy2yvdaFEGR21wuEFsIC3vF1/0O
tcufRcBDeWbiPmg4JwLYKg612LBflQjO/33do5e/wqZGgChzNmaWez5UHrGKr5hCf+IHg4/ZXdSl
rquJUeGZGeimAoW4PBPONNMirfk0ZUlx0adRQqMcqEU+XhwrNQMCQDgyzhpvfny7X6n2X1u7rRfK
TH25ts4SPQ1j31GL/hXA31dt+FUQidJYreUMAKpdmrhccc2EZJOi1s+sjvoLelegs3PInzxWYRiS
qQxhg+8G5uDv13Cg72fBeR97NvJZ7Gtr/3LQxR2mDdMHbFukXr9oGf+KpL48o9I7OQjnATX1Yt5n
vT6U2KkHFGLJ4cbRWzwtRwRSr0Lsp147bU/O4DdMaHPs8fuGd7n/C5vPe7pzrMNOP4x5ex27hHzH
7CMXzrgGnIA0RLmEX6E4dPTC/SQ/2tGXStrSEMtoa5OBR5NYcJHhANi9QCZKgltPTcgQgiF4Jbyb
uwFVvaidE61oxg1RleEEP48LwxzVA27vLaYsQEQ+UCRv5ka13bL4FBdnoimSG9myZ4oeZUmurqXt
Qj5++2pAiFA7ZR0pM2me3kzNzVFFB35ACIw9IiSNUJzXu2ftiSTDr9+ydS3SPnuE7gjMsZriRufc
hwb65bDnrGpRUEmUiyk4LCevbLevXHvn1PB/GGDE0jHOqkZ+oRqqZsmIjCR9i1fjfevIeMGTWBRI
8wc+f23FlzEdwvZdletBIpYJUUy8RUzYQtpwZ7Pdz6MVIElVjdpyG7j+MgRAyNW3JuFYLzbzHr0A
jQfWwoytk6DDu8cFxazEYHFwyG141lQXk3ELwgnW9Ch8v6dDw7IOmN7ti30PWh6eLv1Mh0aBWA7L
Gf1PP6zkpr5Y5Abf9lXlzpL0fwdG8b08UWJucX4AM46b5NF8tqVFUtJuwBRs+6wgK9y0xJe2q+g7
46Qlx4VoeggBPg2KzG42lMwc+hzeVv3hIlL25F2t9V44lIUHIt+wEvk6pk9wyeNXlkNGiikTbL8Q
3y+j89BW5kEoA9iQUxRhm14v232ljehWd4lclnyiy0XISP28raHEvfTTW5iyOq9UmPx0aT/EgN3f
kbJZuwZUR3lk37nWsRo+XUdVJMiMTD0TZNJMJgdO8DbOMucqtu2FZf5ZiRqaSzmil4z4fc/4hG11
lPFX5TyQxgU+etV89vAmdXdQa0DF+J0nvIZ3IBNbq5KBGF6GYX+Nv96dzUCYhNE++sThGFlbnrj2
pSqINDquepAVoxzIHxWzdpaTPlhoCQPCBA6UHJBZdTLEHelHw6+ekIQrYCAa/GsEJs4ivEMhyPTz
iNZuReVmpYyUjBjkm5yqSdlgYcVxQvn+anvSFtehnJZdrEjsAmajEANXl/sA9n1nnbkPxa++02mH
8gu0UWhpwXhvbCOeQA3iV2v23GlC2pwOe4QWIOd63UgYBcJRpJcY2lEdQavhUS1lsUCbpjjU8aWe
4DJJGmh/X8zQFBmSeZnDARgAQ1UFgVybL643SQ4Wq91ign4sWX4v0fEOoHhOHuomIMpqkqkSN6ls
flqdWb6TKS4WvAJHmj7BG/GeVjNtLt7l25Yrfwm1ZRYGNi3p/hG4ZI8gezWmBN/MriTLfLqMI3o0
EAi77WwzOf2fnVGEw7ngaijfXGXad1jsP82J2w8l8ZcROmpCdwWmvmXf5H3CpJCphygTz8KCxlNc
zJ3KWYWZg7WHvUgDL98tPonvqNb0nv/DQ6irBdIIsW8yNZMD2ozLuoQas8YBg/bb+jtFwN1HkKLT
ds+DM6Aq6DxKuqww5T4O/MFyj1TAflmp0OwIHIT98vgVQnCidBIrpvMysouhZVsEj+i/HA0TUGAk
fi0o83az/oYRCA4f6Ro8Zc1yE/SRLdD2qYNk2EQd/zWK5t+FrR3HU5+KfjYeAOY5/TFxEIQgxNJT
JSgX6iYAbIW6682Zyh7YfJjCHU/mlZ7Zw9zLt5cZ96YiC0iSTosTvihKw9yzPS+lv7gPcixtVqtp
aiY1u/bU437uQB9K+CvKycv2qW6DSMtqOPc0s8sAye5clV54DP2bH+PI4+PPxmTyQO8/bsYQpDYe
RbD11kNWMsGFvjnLGPCcHSAdgD/1xkg9FDw5ONNscWtrEK55wEJp4ciBo4epbB6bNAe7VpGGCEYl
0pFOnrwrVFCbzGUUO8iwsdQpzBVR7FLp3XkbzktVM/QJY8uwlLv+usBaz1Xhnff2kABRa2iKZHLT
XX9WhAeNrpqnqEuj92AqZrNUIzrYF9XTWJK0RWupCawvGz+fKxkKwEbPzJpxPa4QuCU6NWmmCTjC
tsG1Ap1gonsp0bxmXCNuIu7Spq6zSdspz/7kFsw++cuxcl6qPi2Ewc+3LVWulMwV8d5AGR+SeS66
ItzaZUiBZgp4i1IPZQ4aKdSXy0CpQAUiMO42VndEHXysspVxoyC7fZ+rvgV7va1Knf84G4uS9Eat
2Dp+PVUHjjlE3fyk9NkZNuOf03RzD9tJEX2k0y1sk3H35E4yokN+qvn7ilIfTekjD81nkBOhqtm7
KS9IdF5tEaYxE8+xp9IE2XkOZtN7KUuFem1eOaY+M9gErAKs/Be1eqBaqnL2ldyYOMW2ppxrMUdJ
SwSWtDvf4Gf4W2BgbLIXVL7TV60eA/fljiX6QVe4eJND6xih265EbT+ZHyiZLDVSUX4pgy6f3+Tw
4fT+Au5ZTjv9llx7HlSbAtJ/PU7aKbfTPmMVb2clYSl5sxxLZxOgDZg39+WwoL5paPF9R+CLZnu5
mN/HRf7jFBa5MVZ5Hjl7B0v4P5xemxLW+JMBG30N+8Ev/beuCV9H7FwgJvLlVEqpAAlCz+0YeKDk
WpsaQJg1ypYf4FNGGKlCKg6McOyd4SOFPm5bg50TnnmeeijHWBYhpBI14pZ9rn2xjfED7cyBlku5
RxBh9csNaUIe2w+iPa3m84Mxxm4fMHcj9R3BsEVdDZqP2x8d5NLuIXID13ZiD4VWQ7pgHPlzejOF
P5H5jB4gMwWm4i0ojBoA98B+JX1uPkRUzAcbh5gpFnl3FSHfOiGaRg7wZtJuIc5g0LHhC+UV8fPA
sXeAK1VruNtfRHbAyCgo+s7LQ0sLE9X2ne0fOf82HIKvQJ2evpxKcGTo0GlS0WZKdp0Ypw2iaGkY
+jyM1jzs7JH+7dheFUT2fq43tZaksQsoWswCs7mdsu0/zID//8LVSyhkQnAVB5pj6hpDQXNqM10x
gH6aPiLdKQpph00LNADl8opDq4jG9hKTOV+qRuibB35BhsHuYfRD7MF9kfp8n2jZu9MWzN4iYXKP
xEneT59rOtzavWfnK7ZJckEZVZ/DiwUEne1Fp0h06hHaRbVqgyp8YpEMQS6Rp6aRjWKYrKRboTjZ
o9/smm56XgIkZfzGw60g/zZPD5VZlP2qLx3qDzMEEpNHlAvc09BczWu3qMIylt7joYb9FX24CtNq
BfbkMAODUV0sBrG/nSyEu+++3gf/g9M9X6DrrqaG2JkIhah8UY12eNHUZudiVaERjNckJa4Frc1G
dISzqpz59DsXOoznsJKGJ0NQnFqrR0bOIsWVt0qiE0MTQ35uaJNE1L8ZWFZoABGmndDJBbYPDuvD
YdtaBgNnYA3KDV7S5cJ1dWuOpe8dSTZZrkdYGDGVxHOeUOr8M+Bh2sVM391IeeARFKTfH+ZNEtb4
jovBcN3BgLRpnBis7vr6aCR2Yhimu1l7DFmjVStdaVSs7C5Zb2VTgDYzUAiH/tYKo05CTH5yVWyc
u7CMXM7U4KJJ2BInQ5tbNoMm7BawjIVbWehf08nKyGqZlHjAdt0k47MRoBr2Iuqz7M+5TLb2XxfM
L9ktjVm/zmtm6uBQAOcTlipbaMtIaS4Ek5JWujb2jaNQpF9xtBOWPqGXQpZ99sE0iLogCnumvFxY
dXzZrNccIihoCoz2MvkbBYoLDKKzD6inRLIxspBzUzxOoerfX+4ARHo/s/s49RCmxqUSYaqTrrTD
9Dq28/qAO+079+QLfdFHhH5vENCyz4ZfV1AMfYRvtaxzhKvvqepT7s7lRqt/N4dnXl/gA4O7aNSA
8uxXjV6Zd4lwCbYb4sBa8+b2jrZObK5vOS88dVRFHGc+xdw0Nmx80Sh5g62Ul3LTA3NhQqWVRT9/
nnu2Ah/3YXV/i46PAoE4vKyIkEINaLtdDEvZSu9NaKB2tSAM94/NjL0P6kPPz0YwQ1/HHivc60mI
FZe3tI0VgGognFehRO4/HNSusAEs3CM4WG3awvSnzWvGcQsVGrqrZ2Amlwl/bady/y57w5hwnt7L
PwHbHRhryigce0bp2jVV8+zqnNBnVZTACsqmDALBZxTYTFNEHziX8JpfM96nRcBk/goRF2+WxpLe
frr8EwMg6+V2y19HmAz8wqi2rSKjroT2VAf9H+M6Plv1vgfwbaZCDZkzoXBDtJMXa0UfL+GaV9Rk
hv1Kj4Sjrka0V7aKCoMYLU8BO7cIzE2oKvRJwlUivgxqYY+F+XYPYIhBm/OxeAW1Nwl+/b61TCb8
0QsiqfpUZl8P+J2YOolmllDRPHdPT3zkhCWZniHZsAGo+8NXJawvz3fW1yEUvfsrF4O0KBA7beJ0
2gNkJkwaBeu4n9DFCu/ug61g9te5Pu6mTHKqdG8Mglmd4ED1SvfVNTwwXG+rPdtHoaEiP2sy9iAU
O0Ny8ToeOhq7TtkOXsUiLGJVJVmw2h76CfcfOmH3UGRgdBcl28wPee9BR21W5NwjKe2nh4/Mq4lV
lkOXEIRzNaMwMMfoyXsiXz+P+4ltA5ah978UAERh/eLHh367swOYoNwOEQUPMQUOYAdkPPBlU1MS
TDZ/IMm3VPHv7n+b1lYWHx2qdYLqASTfGr+oeYygJI0p1Txe4GWhTgHgofwDBstNSUzCzguq8GBw
dtu+C+6wp+1F8kD9c7XTc8hTmwwU6aXhZzJQULGIQgOtymq1CxmbHFT0L5whOTck6tM6GxRcVuKl
+IBizCCGSMbJdEobGeFWR3oWBUIq6FVZ+uZAVjM8DBkxVU0W/TRXV1toSeuBW7eBl6DNLnma56SD
NlSE0R/R4bU8MetiKUYqOFBpBsEGmrL4AKI3bCzi+lcYj23BnXr4TvliYW36d3xkq7pHtEsMMXG5
ORfXZyzk6QiLNW9TRvuhDBFUuefpbEPNEmQ+OOccKVoVYJRYS+2JegMD0LMtNkwgQ8jb7BqcTsrH
HdOVWTk9zrf27aoR+02P39cRgPYvE7XDMr1VL73Jdp+QgfvJwr3Y6ksnIDcUO6Y+2eY2vEbtFedy
oMNo4nrV29EgMC1eWx019Iq0UupLNaMO9ucJN60dDh5u2c1yqpOHnvEuttegnm/helyI0tyGgQCC
oOU+bYUvOgnYxMMP6LOz/XafgUT9yJ3GAoNsN/EkPL5DddfboCfe0KTuTbJVvnKK/ox+qtJpke8o
f7ITxxKyiFmG9Jyut09K9Y4IZZLdybnbZk2uhmb2KlFkGaxYDjWGU3NdpgXa8tQdh6OqFs9VgFpQ
nwdWI2Qu8rKfetvdiT0QO8pfhzHUg0cznXmdiioxiOjOEl4ZmJvqSNCdf+rpmyWBhgZSFkLERXlQ
3ZsGMNqZeJW7KXbmWkNe80LmZtdYkfZpfFVJu0lIhLtkSracfALeaoMbbpoT+M0GsftE4ZrwJtE0
cZYk5iwvbp8djfkpVb4BwnKgxRpR+5hqDqOGVIwgW1K4Nz9Y+t/ybVNCb/clVXx8YDuHxEFV/pEZ
hsVpC+lXCEesmMT+jFTVEfGd3O4FJjuv401QFgQWHBPEKHLBgWJmfphHNLl0r1gF3aqMGRABOAA0
QVBC93P0dtoLLvhz/ynPnyrnFzXiku7mRNrdRNC5Amr4zPco0CMm80ZZQSuVPPMkx/o3BEp6fkCY
8rj/c0Lm8hAbppQnSNDqsIZOOjxHwBVd/j9VUxZDzdjHu+LiUqXxwxVFjLLACo0YYEfQjvd7NGSr
VCEXD6+ayuJe/0C6fvi11006k13kmW77j5pPGWrvgSp+G4+nE2WADUA3lKhDllwZEE9k7vM2ILZS
cEvKsBrkB3lVBsBDaoYwfpZp0SP+NUjA9C8uQpudyRIbwtUzaAqTQ86IV9fexA4rXDbV/eGV7zpN
l+LIBvvLvwPzD3CJ9UfjEc6BEWu2suMmThS4yujuFaWfRu9ipRlnLIy/JRJIdMyXuE0k7Ia+cROp
ly08PCda/xr10NnrEEFDo2VSl+rxP6AzsTMpMop4/3/5gt4uSj2S2LtIZl1l5zyVQU4zh7Ho5uYi
pBoD5J2elfXSmqm6pEZGKbgzU2kmRoG0IlQgDdnNzonM0orgCoTqV/R3/KhAJEtXf8pSNIG8yoWQ
A8l+Cv9/JEN5ucc4W4YK6QSZJbMFmQjYNMi+1lO4j7i2FHbmBTY/F/0Ru/+s1U43btUCQUdh9ZBU
8a/UCnvBaRz30f/UdlRGHv0wOngG3py6Ce9JyfOGQKGwEl9gWdQkSLhtuBIC0qMqixi4Wjg9CyQU
3GP5PV+4mdW+VfbXBFm+a/aHL+V1sKy5dWYOcAwjElclW2hnJQIM1ZK2gOqQnYWg1UGFSUasKuTh
46LUnq2kflsNpYP+i68wqA9xhwFIkwpxLhQbxPtsFIoiO3UNE/bJSoAcgU5NWrvJQWz5LUzy13UK
mHz0RaiftrM9cciHbwMZMZzScdJ7eHsKqRUILIakvoHGQ9kWt5uJButeG8KK/ZyTyy4UOjbrsL7V
EdD/QXaWR09DtiMSF75nD5OKJuRH64i03624tEiPN/6tmeF9zYxby3jXeKnjsdE37tcc6htcuaR1
i2vEMaBILPqXSK+jfFBdoF+Sojl1hQUq6Jx3O5VVEDCk8KgkBQfFW6BzHX7lzXb8mMuhhEjz7k5Y
IauwvKBUeH7zzFWJYJ3i196phJzfbV0C99YwmFVo9zBBFgZvYx9s+m7mHDzgQTN/sey9E3+vikhs
V6SHcC0O4S+IAlr/F3FgjNBbpFTMxKspTUbnXZpsvuphY8/7N4qESB7ax8JGnZOygqnfcsJBGHGA
wyUHN7czSW4MHLBI+UXUwg8WDRkZE3tUJ5SNmx7veFcc8dY/t1blpW2S8WcBiL4qH6Zd01AUk51Z
egfKqWp8XmFannK26V1fqzM7upZuIRIDo53YhAN3FgKREH8JNE4V+P2FtV3ml8En0QSXIQtADpkh
lsZ8gru+dpKY8H6UhDnY6uLuCMkHVTQoL1ptxnNRtPclbLiaQ0LiJxCUMaXJqp0jU/k2+azL2rZ3
An4n/pJu+dCeYQQ7MqwjZY1Bc8nBpTyeBKcVid1IrP8afump5LnF1+a5ux63shl6QfMOV7+WIX13
L16WcIljGIhFIazaTZb36UfnoHB16gfASbl3JNqXskjHxCeA9Gag16W5K5DCrcSVdbQUcpf5TrgO
AeRxiKEN7N04AQ4lfVinUh4+1pazUwuooWk6fJar53jUo9rrv/AAL/n2+B9PLbOmhtUH1s6cfrjM
pFJpi9cuxqNUWC/IOWNrx/h0VYAGtNTUfN2AJWUEbKwKz3FBzIW0trsLkZ/q+vbYbyp426i8uXNk
bpOhy4YWEVrzlD1IS2YCZsENS7ishz7f+O14XM85k98w7X9yof9bn7Sab9dIXuWtBIZTAzX/cUDP
bNzJQA0AHImUqJFFZRLBQlV2lTqrMQgm/ilqa6JNl8xNkU9202wIVO1jfovva2FD4hvUWKooGQTq
abEbi5C7W2vZurKdQnj3GfCvc+TbQ1trOkt6IYffVKIoJkOwmSIbr/FpQZ7IP03fW/82j/wO9646
GItpc6qDXNrE2NjVHJNv2dPy5HAXkdP5Kbd1Iwu05DnKylEhFRsyCnIjjkYbijpCFPrHlHClamkp
QKY8BRz9nKmoNVh5i8wFvALDUDJ/wdawH/l0w3drXH6y9Un2i62FZEahKI1c+ldpbeFA0/S5NBTO
ra5CiQ44AnqpKg05UL4SE/r5gJ3iR+xyz9BmfqY9VtoA25mytUMN+sCcCJQOp3HZufzOfhr1KL+j
B7/fCSbkb9mVFMYRuLXzqyZyZ01I5q1yRq5tu/juw6+/J9k3gvlCPFcBJSDOWHG3qM7YP/Izr/1a
hyKQB9ZltZh6vhKNZHzz5gFHe07FGq6EZhHNIWKvWCF/xN+Yei/gV2GV94c6GLRLjBU4zqTamFmw
9AR40Kp2V8dg6SH+abKeBveGv2dRljkwbYxipXj2RKBIR2X0oO6jaIIfgAAKV249rLWo40U0Dzh+
Klor5TpOPCX+zNFq0LaGxI2f/J0eScTy7RUEcdvdjK03wyWuPOteMBCFPVHGz5S3WMEIR9nWLRk1
UZD4HSdHDFJ2NQBIknCDsIWhazBHNWyYCaI8A+hfAd636fpuvFeFMZi23OUe7pvwSpLYIet8jZVZ
AcQP6p70l3J2OztAJ3q2Kz/ABhdeV6QLtCBQYQ/n2NJm4ebW2LR4mrJr/LS75A1o6SfzwO8TN3zX
yDKJNoFSsZtcNRJwvCqz9q7gmWj/6a5oVfm5w66my/JhtDRUYCfZDZXJ8WrjCTcNSM5ofYqoJSBe
BDs1lPLTXsYPBS6sDsJpvCtaHB2xOLt+5hQ6+fhoVXaAse0HNVColHMfQH2DfkLmLcF5ddoxJxut
SGvADD2SylTO5pqBse6oUa2psC9HQg1hRLVWvHX5z1MVVOVsvCWbhJXEs0+iTJik7Pqx4mj1dKbB
8PnIrzxfnwjYw+YSTKeVEdtMODv85hDUrirvCxL8hemktN2M1j28cguNARnKkYDb3wy24bObPevN
miP1BVyCafW05tpxJxeZrhtxoOWe4586+AYKjGWnCo3iWb1SmXa1quPQQICZWNqzPcNttvvalcqW
9UTTPkkH8DQqN6Am3EHDHlu46I2faCUm9VVQtSOajOguumuI1+Iz4jNHHgrPBxRgFjvNciedygL2
DAGQmofrnvykDJrnHeOgsCOnjsIVdCPRK52IxUCnrmY/prLmgIKttPEZ2BbGP4uMl08Y2aFWHK02
dM/pOO8AhWoQajqnJVepxu0DMFo8BxgJhuuXPfERGPLJQQ/jwLyCzNjzGIVNiwDZt2Pmn4QMgr7N
d4GNpWsKt908aBvNmorzd3D1DlopzYL6FXPS24HV+k9AVfLKuv2lNd5ij6YoyK8Vg9zaEi0xIbbs
iq2grf2OHwvR1ttlegFkiBfGSkcT0l26nWVhg+i6WqP48NwapQm4jAncuHHX4N0hPP8qnQCGrc00
ATyCvc5tne+3G2jNY8GqduA/i0LY+tRmizc3PDPhMs1NNiALkEkblip2PSLBN1UrBeswZiA6JJdZ
S3RreTWaiAkP/mRPbp4ofZTYvGXocTzC2WUtQiJTg9sIU53GyM7B6e9b0Kz0q+3oHfrWUzTkpCPU
7+Op9cYpqvHlb6Kwrc35uzXwj1HuZr2Lisi5zLnrGCIcPnhV6Bg0Qe0/JLaP88Bk67ACDuHlVBBW
CwafBaSlbtpMCdwc7WBTCMlNoQBlMeAoUG44ylw0pRz7P6ukl2XjpYFPQhV7oNc5e48a/T7gOeEH
JIvc7+apR4Ha5AnjoWwc2jgW4Vt0oJCheRC4XuQbvNzJQRz3qLEoOAyii714a4/5L6zHLI8c3GNF
GyAEWtB7ncGfrow5GkRSjj4QQLlFSfnQR+6Yz1lEVmlc70zxFNPle74zgO/em6X42UmUZHPsV6la
nfjtaclNZH9yjZpUG45XNXB7xlriM4FqQbxTHIUTQkZ9grRGbum4supUq2x4Umu08QIk3L10BUCK
rlPl+z+LQ3rtraaF7s5bTUqR2dkvuIQnS1BBBsu9Whw7zOVjmlxNrDYSMKSR5tRhYnMw1WQtN0zE
T3PKaXDFUM7PETPcNsH5jd55uL1kcXbWsrs3COSaB+D+6mDbhsP5vxDWJnJA4BX0juZCsMeigvmP
1qPklBmX9KywdD7jNIKCZr+TBWhjgB+wxje4ChgSx+FJYyosr0rINBffnMy8SyEr6ajz3U2CIEeS
KrFcdqE1hHQC1wALWUigCUZDVGw7qLQ3ct/I5anhuq8zqshjeMx6T6JFM+NCG+OiVeCjEfQu6D8J
7o5XAtFtXsOapAZmA4vUWE5xL5Ea1abyJhKI7MOSRK1hgkj0777m4B4CAjFYJPAJKOh22nGFZIXk
zKjBUKbGhlqxwgv1dnZlmvFtQIjIVbBi1at1L5Hmcl5eJu/bETUb15xhqJvSrb8N7Cfa5dD79zpF
tILZvrHDJcChzRu5vM6H+x16AU2fmNWXsuoXZ+m+ieIPeY7siBnHo3kG7aY3hiz440CQwSy8Pwjm
DHzq7boJrY7DXW2WclUDkFDjf9zr07HD0d27d2iuOdqAHXnVGNab0LPWSCXl7SpcIpyD7v4i8TmA
79vmzZ+++LqGft/nmJaZiZI524PSGZ9nexgCvznXgGLHFvEQ+Ss+TUVzZVxsAC7KCQ+IR9+vHsvK
HUsZnRWKgw9tEtAi8muoDxjfmMtMDcmPA2h+AftZbVulGobN8hRJBZrFuowLGZs/2UAQxy5rovK3
TLMxQGKHI3msmZMj4Uyi2rqLioS4muyvk1q9HTO09kre4oJqny1AzNELtPiYH2W4EoKIshJy/z1x
G4ilFxItDmEdSfN8H3B2xGyAfGCPZcwPAhR+PKrmtRhNt7IMiorqKIW1BcuWKcT/jOvNdCGLQ5x/
7nRpjkCxwK0F2rsLkBdpAx2b1gN/y1QPYaq6oVqdZC9YywOEZrijrTHvPhuBW4bqRIMhiGsd6qg8
IZ6Datle0GFP6KNkMtgB6d6Z45dAOpYvny3HOZaKFH9UFppvFlxkZETkxJGhXFGZ27TzdNV0YwV2
XRlunXA6TQKl3t0cActOKO9LjJfqGjy5ANynjKxoYjMeJwlBqERFxxfN+cPZ2fKrDS3ivM4rNjXz
N9RpA6ZlPZtwaoWZRS8KgXO/DofJh1B0yRLvDu8bJ2Jdxss3hMKrZEDnuMYonPCQAyl0uAGTnNLl
4NQdqke/04MIb9qGkumspzhl0XLpIPjn85PrJoVyK9DKuJZtqtu6t4bfjd4+zKrahxVQvxHUo6SM
Uq3y0zsMUnMLOmJUZp6FTQdPuJ3jN+Xsy3RzjhAbRViuA+oQ3r8sG7vvY1sCnSi+fLLlRUN8FXXG
NAj5KEuwo9q2ggzne1cjJ0nDGl20fvFtJEmHkiozAoBrSMnvfIWOWGGTNHP9cLYBVpTJvmO64IKZ
QSTCSgcCY90ozM+i+zar664YdEwYph/zF9rGnL6qh7b2hJO+CAvhz/beJo2V7ePhwbuMtYkx7CaY
yt8tLTiReCDA1YPCWDpXccH39oH3WGDSuvyC+U5XUtDmDMcUyz0QEdTkczYgIvoLLz6kSbpyarjS
8ZbnhuO1NEMw/NKEl/IY/By7t53O5x6PgltFk9r/6vp7G61EpkEL4VNAhPZZK2KAD7kadnXQfrKv
2FjEdsAlwB7dOPUjt/5kjKNI1PNZ0ZRtvGckx82VTGELzr3xNYrnaGO5DJfWiPHIap51p+Ckk03+
SoFxC0wKHzORj1YGACSnfpx2BppqbMUx5fpbGFRRo8UwRWYG/1vbu832iHBXwtXUeIZ1F2mzI0Ux
X7H0reOlNc38s0+i+KSLvM0HZZ1HeyXrB8Lk2SLV+2ug06MIwH5LC6ZKDGn0/bIT6J8sLZsq778O
gjhUzDB95n4Xnd6Jt1OcpjmhNQFwjxNsmJHD3MvA6n2zDDoZfa8uSVe8jUZ1/YUNs8ky7z+C/Dpk
cIMdyk0EBaGRxJn9impcu9rIHH/9DTDP8qqAmEcNusDCDmjVhA4HXZ6AmrYcNek5vFxdpkAtR+kk
0NMJaeRsLYHREp03kb/Vdu5ayBqzxzrfYI/vqUP6NZMlheHT7tamuXD1TEseoExSVDZKYlk25ws0
CN+Vrx2/DBfgP2e7j8zVVi0ToxCRkk261NfXbHxXLehI6yRTi8icSpP5t+e7nCZ5SzJROYpzzaDk
x5KxgLNN/z4M3hVRULdURFLwC7Ift1yn6y5ba/55iWHTlG6u/7iqZ3Xx0Km3gBRY26u75pi8R8ew
m0dWjykcn4q/bkb2iAnEBpc7vYn0R4YXOKj+Yi9NwJj9+EdYAKEB089TFW5t2akBM13vS9qb/VWd
QZF3o5WHHpE9UQIAiPwd1C4JsG7roZcNRUC9e+KAUIBmym2fgCuk2+/oDvU/r2EeY6p0uE0WlKn3
CIrgoa4SyMvt9M9kgMgYPmNT75V1giGftUMiQJr79kLbnPcH/vJxi19ow/mTFr1XyT2F8K45K1n6
BOfnJ03NJnC+dpYoA2x+pqusIlleNlE7kMNd+pXXweCHdxOfdzbVx5ZL1ywCqvF2AVqEZt3QSXhA
LoeNv36JoppuG8ei6XZXwMjtVnHc42h67IaTWdxMd2y1HFU3hDJU52l35r9eBYdhqTL5SJtRg8Ly
Fnfdx0yGWIdNpKaguKinoy8wtiNbK7jShjTnLkypaGNcH+xRX+H7rYO70CXsmeR+p3xVb2NQ2PAP
EyZN4/K5X+JDZEDgN6qsGwbAdOtUHza1KgBkeKlAYApC0fxmnbPMisAxVsnD+LTbfQeWaqAEPFTc
2ZLrsHkvTf2h6AJ3M+gwiaXOYP/ZGEZ+XOK3KnKEgf0IV0V/CzCfRLto55rhy22xL2V3tyAXlcFH
X2raVj3gUWveGJDJyGgdYgulTRruIJ4kDTDnFglTh4qvppis9AOMWf6Ed4FLmHhQECH2PTSBowEe
1XlvilY2M+5IFEB6XX1KQQGVpbzvXYbHtu4HP0Wx+XQaH5F/G81SNsBsdy79EQfXOP0KN/kHwCdq
waP5vC8UlIl5/ssqfBpzHPMXi3qCbEJzuEiTGHS2sQA4/yc4M5BS0YrbYF9QIYXV9OQt+LdIjL8N
LNqiOsKuvu82lRk4lf5ZucB+OZdnTge1Q1yVS4kRMSfnAT9elj9a2X1h4yof1ef+Z1SwfbyXf3Wr
DsjevIv25HtorwNXSvbcTlhEJoDd5WYJAOzkL2mer117ssq3H1ELKYYaDwL5MmOzU6OGN5CHVRd6
huCDBMeeNvB3Ig+eEclWEjag3MVWmMapseYESwh3ATxRfsir+/WOzF/nUDuM8NlUHJCvFTwQAmXG
xQP6TDQgYC4vCp3m6gbyzo469BU7pA5bNS8YfgqaBtTt7ekgGyPFbrrBrjG1HNKas5an/BuZOPNO
zkdI48gyiahI+14Geecme9M3psXuNMTuCJMNHSQLDDrmM2LWzfUYgmgGBF4aqPjC+7TNppBecZ6k
u1biJkml7M3/0mLhOCENqEk1jDk4QkD057QLyAF47rWeR3VvSpeIvDN2UcBEFJ8TM4qdP4GhDG4s
CkUduDv4VyEUZLOjeVysI7D0Qiy20bW0BQM4ELjA6w2H1YufnfLyEPQwjUbOx0yhYerakcC5TTWZ
Orw26PYs9pulEy4FHUJrJi0mwwA7Kbub+pDKqrvvdHPLxnHq5RoF4lT0/yzdkhZm3PiXcm+JByYK
2qxFZwoFIfX48Kw2L9aAN8alfQDq6mPqTk93NvjSq1qIMrMhHMrWmSFETSPNNlE6oKLj+nCdBJGq
493vko1V3FGafZ+K3wvGmvO04widwyNeAYprHq4MbYLHtOyoyC4FJoeMlR+Lgr48WkydsXAdv+Gr
CDnBKzxLg9jCCb/9ZX2lgpDA35BRAnE469C3zmYL7i36YjQI/s6ExOWJ0wUDnhdWoSp3y/dhwOZd
QPx12nfyRCF2fR0uCcq8N3VLqtNKpB7zdaT9exjFFuleOGmpZ7I5GO5brk2ocf6fkL5d5bMQoz7B
Xpjm95fIhPrc8U7ctSAtsn62O/OAeMyS44m2PkncGYFMhP754DiVyN9/gZy1BMzopdXpy5CTVyac
7tuwvcaQ4/01q/LN9bQQC5MwvoWujYi9E3yJRFULASdBEQHyOxmgz3u3AWQJMVRuC0JdQtPHTGTL
XUgtM0YnuvHRUVILRWUkXqE80lVUkXJx8YAUiRlap77APf9ajpTvcNTEBXpdy6MAua+UnINusqA5
TQvGgGgAuotFWjHr1qqgQBdewfZECx7YI4qRxgob0Y6cf6uRXVO8E7Cbju7E4Ue+RIaJFYR0++jT
Zpfqw7qJ/97aqxZr+IAn52EXA9edb4TUcxcAVkC2oaerM9oWhc1FXJ9q5Q1V3Pp9rgr003JMvxcu
iDNwyZ59m/gJAGyEl7ZlWMaUDryhdN1fRB0b02RWREex6ymeTTD0nxcH2dfPt+UIP3q95JteMc2I
XSbtbs/vkFUaa6gyhH894ewnk9E1npO+/nXYxbgjAEaKyLffvbJCOpv5JOIkOZ0M84HHSO0qbvvN
Zcb1NGfvWviAl/qi1WDrBwxzaF0ENKJK52U1RHvdmWy/kB8MQKZhTsOhTxkmGO4iN9nH9Lwme+25
odhqxGzY/YBVSuwhw+E0CpZk31QzrwyRFNAWr4ZhVjCOEEck9EzaPOvjIDK0JRFZ436+FTOgzdpx
xvONOuFnQnt0SI76kE+qS9m+B3NnBKx0sHJc5mchOmYk0GYeWGcpA+ZRkbD9XRmNjBVGpLG2P2Es
2IJgmpIKzLEPuzfBiGyfuEQOpFo3/5yzJw8rIEtCpXLLVBUzUN6YQT5KMWtXraCU7oWtr4qsn59C
JCiYmAlPOkCp/5MvGCYLxmX+avh80bgjAx62kOStN77pXlgOV7Ww60ZyYSxJ3yxAlFrz7Fnt7YTo
Kmg3JmtLmjjvRIRwSrbcPPkxzJ4Cz6Te5cPHX8UbwiYyymMMBHX/0bVmoPp2dqAoSQBH7Aqx39hM
wsuky9hxeAvVTEoNpBWOE+k0uOc5gJ3z4yrdbjr/aEaJwQr7+p1RRoMSzFHbAtzWotnLWZ5LaRh5
Qs7sv4DuC+P2kdBRJkwPh3Pe5wxOtqgIGpfba2eMfCteQ8uX/8BBemzkmGU4nXJzQNtN02UweFuI
Zzz0vO6633GeGIjtBl1ujwdEtK1EkX4wtJcpQTamOb20A3n18b3TVP3BAXYAaEE9kjcvOI7RjNYE
JAEFgk8K+MYWoQ18n9LXnHXWSE/gNhaL54DkFcVWpiPmbPCStqU7QpLVynsffao9euFJpRq/AGUT
VYhPlFXbU21UHAmVzOxLh/lqRrHwsxtTg9iiTXoXTLrQqsqfW2LkRL+w/Hs3fG9s4uGYvjUG9EsX
ld8EorWPrnVIlHKXxXZ2t2wzGu36hgVOXkvX8JA5cwvkqv9aWlmHy00I1KqSjr1LRIQw4P0zSpHn
eYGXBR4y93Z2RfTehRdqhdDO2RJfzIlcxxWvbu7AeIlubTimPIlUIOGjZ+Jd+tvuwkzOxoHRiECj
LPyE0ayxAjSBxxEx6PC9z/qk7tXtKTZBdvWuX9qGUMiAVdELhhK4D0s4VJFGbdfi0Ds2gwvX6Lmk
yOyMR7fSkFPm4Hl+yA7sudXICG8y3q+kNu3FWg4R8JBzZDaLEn4hsClZdrLopvDz4Rfi5rOjLk5Z
vb1a3kGpd3zo27a3H2FhGWc39DIr+FRGkJTUqAsfsNXsVVPxw2krmvOqOf8I2/SjyIYv1U4/TsNu
aLzqcUa/s/zEYhgUTdithx6ESyMnXAYMmdfixL/+1mLlRSIwvUPheNZZ2EXtRNlso3o65vx8Qmda
Ky/Mg25+oCI8P8ZE8Nhbq4AlAQx5OL2XyfBAfaRBt/K/W5aYJpWOTGRCNHMK5Gx8wJkj/BDUO4hP
gRAxELaIYyWxUuEq90pqsnvVyE5Ncbl+/peqqURcHGq6OzP073tC0txjh+kcjIVexPc3OjmMCpob
n4nAH1ufrUL63aAxZD4WfbeqNXZpOo1D2YclBtsVs4JwggISv/87qfozBOexu2D4luIRvbxsXiqw
F+yaqJEaUgT+VsVinVXCzA1ZpkFNn9lT1H2BJDfB2n3Swp5dgF1uhpG/55GPDnN8suX/6BfF9LAq
Ochgwxi3nfmEVMWANg/WkAB5yDgshP0QWZkNIyWnxAZAqNqfZuxHeCBDRaySDGqF5NqPHYL4ULe5
8EVKnEFcCgpBvyzcf2/SU7DJegF0G3q9c5vYGEaFR4in/sOa1TnCB20T/qQ67/eV64G5XMnQhZNA
yh9fn6w44ear3lk/DFO9P91BmVeLLlXgQyhb37xD0yjw9N91Gk1ygRDMQXLuHqWmrL3fh/FB5KCU
2+ofL8Lmrw7WRq8KOiAhssvJDPfhz6JPW77+y0jnx4VwafexlgpknodyVH5cdieruV8hGlzCcL1H
RiAv1YD66vEjbxF0hRQEPmevSKxxuGDJgaT39prUAnLWRmYl3I5H+CSOHU6BpxFPm78v7rFiDOkw
fSqFB4ykJyWSSX0elfySN5vsAV+jAXkTJvic0nmi1zruQOVQuVpTu+oQmHQXZcYbNOLgPSBcYQAU
Fpq/dd4+yTCqUVqsAZOdxPYVR0lEEG5DQcPnTHR+l6Ni8bu1xD4OJMSncjnamDtejwrTgjHGoTbd
1U8IUy/T98zAaN1ypTPytDwGvu+bc1X8fb3F/VzUJrCWrVQOvqSUiqqq5SEdoJj/uOtk5y4d5POW
/IFWR1znJZ+2oKmJdx0xW+S/6fKQ0OGRM+5wYK3C0sBw9cz8zuH6WdhMxuXfbQ2uDGSVmIdyGKpi
h7IHWBUUP6GlwA61mAO3Ku4Ke+Vdre2qoRsaAQwteWkfBuI0DlcfTGwwMNQZFht/B3sRHHwUM4jo
MMJCgCoMEB0CgsHx9+Tvuhb+cuYE/brIYjONorCo6Vdg7Rno6BriRK7LRsao7REKM9X/aT+ohTO/
QFYaqZAcnyxFWKaLT0+4K0tvRLiMGlWuzmhkuGNYp8/1Dp31Uo25cGiuxzgwRbUQyisaNE3ahTfq
8vUUAenXyKiDaPxGpN7jYaHO6BPQZeLTDLO/jejd4t7GYPPmzw7apZdZNEgmuOiQRbxwGBxM2b9C
lE8cFIaxP06FvUiPGrjWKa5G9zFIvUedWPFfa9JUxAMi9Z68v67IKbF2QttD8vfjpdu/rNQWg1aO
ziB8VsVKpWr+tax0BkWOYNHp+5gJnzqVyKLD+dj0NecrqbP0OovhZMq7uytWHiuCgCSlkD4DMZk+
l31iBMosCInrj9Rru3Q+SpIPw7mxWCPVhuRynvaoFfGfxN8k1j+Y/oODuUy1Yk+XjMCz9yo55pcw
vnnUdjWa4QnYZOQUm22mBobzQaC14UBWzv5jNrUbVebDFbi8cDaPLYwZJAK1BJI1TVr0KkTkoLkv
PXmiLVeV+tJowWLhNXI2xXR6so2xujS5/F7aj1d05uhyQsyWY4hBWt9E1fOamjcyXFQXhpz3RJIM
py0dlANtAP0mUh6mORmYC3DLfhh01DSwdTzCy/5JRcyQB0tNbINUUAQtt6OSUMbgd6DdeLY5sQgs
5oOuGOmKsJowfGHhuP/k8dFZfye9OyD5z0sMzzOwZP3b0eHNnZl93rmOvnGjlkQL+5MI+0oPwCpu
Q5olr6Fy0CbYiOLFF1mfAGrwH0SkWSyqglqmOT2VuNgDkc1yRbr2nxZOsIRsu0uGRdDiikahmW7Q
wv2Oiz1hFgwVV7xGS8gKQm980+C0HQjcqEkYqChvuC6JZu5X/DkDGwFtVpG7YR83C53oolvGZXPj
OOf4U1xmVysXAdhpqkW61ECmi0T2Va2gsBO0I42UKsqev3uHGOMQ2U+cSt4vfbisbrdo8g+YznTl
kMEhQnOTSy3nRAGfQMmXqQU6Al7uWf+L8PVPP/fCuYswVZCTZLS/PVUNVJWhS0datMgpvxnPZPuU
j3Ke5rtReM2cDT0IZBlhl23XK7bt8pVKfV0HrCODnyip0DLWL8NgkE7HRe1idi5av23EQmwqknkl
NfJ88mz6NkRQVFKMaH+8u0EAOQja0w+mk2XKwRh4LPAv3LIaMmj/K9nr8SWNYVkUSTV1ipioxqri
dlXnpUQnn4lVPc36hqfLjLoj9ei8Y3xbPt+1g/hqm1yK8jndAvvQ+5tX0j+sBc06rYQT3t9xPJkB
xPqCjZfca/zoIbGlScXAmwKxXn+l6GaTmqMAN71QErERy+pSnDT7Z5j/7/8yoIO27yLgwJBaKxye
ETqs8lkbm85+rGN3/1Jpwfz3mYfsm/6mH8DpO113rEDNV8Ty/iuYo7cEkDH7bbp+djfzzVH8h4X7
xDMdoPTwlGEoZOkO/5fWCOpuISn9jXwzrod9pU7tsJqnpiAscx3vDEHk4MaX0Bu5yt4nAQQbHDw7
LCzWFcdyn2t/4aYUZt9Yk6yDwi8zgM1N5rbY/c5wJQ5fQDUYt/An3U9iI1b48Hm9P64MNQYIdc0p
Ooko7O94NydGy+TU5VHc57ImJ1wGWRy+bFL5tcbvLOKGqQ9uU6rb4+PmAO+fbSShqJQqr8hwu8pa
lPid1Q5Z6+tmfP4VWSxUw/Piuu53UW5GOPhRfzNncON39APABzb/vxzKGqxHZje6EqjvXTGqwYos
mrnVaaVqNLksD1vL91L6IKF9tybkYsCBBRTklvxmJkMaG45pLUmDkpjsUSr1HGaXHIbWo/GGpDxD
wd9aru5JOm6GBo+vMcZv3/D9PO6y7JkjDDZoQAMhpUrAT4vp+Hnau7jBNjv9YgLKWQrZL+Z/7Ny8
NLJpMgASZUnjIjnJdI+c2xOUvlPoq+MLU2fLrVVKwxgkncYzDvqBwwZZK4Bh9j868Y0YIbAfd0rD
OaotMtO/AdogLtAWZnzkJS3IXvxpROv4Y5o5gLefnIivkmlY8wn+ogxtfk1ZbeWU6tevVo1ZS+ib
mp3BAwGtacTxJnSE7M7sVbOF3KG4rv0eKBE6MwCGE0ayUhS7t+Ejc/X4rvEX1CmQd4ULD4THIROp
9sOWpN6fsynXAevt7gdp3n3vmOR2rq54GKYgVlk4TB0UXDkR2Y0LRqT/vB/J2/VgTdajpLZvwxHZ
QrXcctdTap8+gDixpCcrE4nCP5/ELb8Nuqo3clY6gvU/hleO2QLoRwa6z0jK9SSHdG2aDKrBnnKW
HpG1XBuuTymWA1iyuKgQD2yBAPvF2VJsFiuKrTanu1S7swg1GvjuayuidfIQxKNsh8BBEwkkWkwt
b6kZkxxwvVI42/jC9BG8zdpOd9ucRCEiJFMHUZj6Gni+ghhpHLYu1VW2WT1vhMBRtxt34btO+CN5
X2ml452IAfMsR3h0iTiNKkM8bNcicMz6s+fvmxCuvetZc3OZZ6zix0QPddAcDnyn1T0ErjP9YD+G
ZkWtM1Ky3pcY42vs1H0O/PU4VrWn2lfy0NC3F80SGLQdYVxwc4s4QWbHnfOJYxtZy6YVbjYWZ/pE
LVi/fZiCpMEgAZV5LlwEHZARkncbhLoUsqg47bvSBQxXzgnKk1WRyViloLTRWcpv//s6n2op9BPw
CB/USkcQ15d5VNKXU5UOJRLPrl+ziviYRyo3sdFJFcfSg0lT0Ba19NHG8pp9qUGXX8+S3vTw1BjI
JF0y3kn0F70g7ZJzY/j1jKIthzbgczup0i882OITAR/MxRBixbJDcQUzINGSVwI0xtWtz+7DRcjm
ImjCRhlFZlA/tsnl1+W4bTJMuhMYz0OHSZLFjiI/fxvoQkZ6Y6PRMXYkzeDBU2HLy6aTnzMpD2Yl
NdEeKWc+YAgfuYidbFh30LLl01i7PyuYmOvUH6UkIxW2Hqeu/f6pl+SmPL6CcZh1wBrzYB/4VhQu
scxlI5/bcpsHL6QT8oqp60bRfDAn9Jskz9NJ2cbwr6wXERXavghaEZj3l/07uLq1S40ZW31AkdB7
hT9RfJslP+mtku4dJHlFbEKThHZm5w6YluKzB2KQR3ZLcYpI2H2HF5cVo1eadWtQsIjMVZn0mZIn
FjmTAqOw6Lyulqh0TPY2L40l3B+a1vsp/DlslFN39jZDuHxc4TX5HsV8BcM5CSrpmRvlMMhMvDmc
I0v55wEVt4DN5C/WtAazWOtSUZ5jGLWz/8BzzJdHEj3LLABVt5QJH76jAhSX7B0DlK7CKxPvugmX
RaumR51U5J9U5Hdk20ejO2dCPuhq/W4UlIK8+8FH7mkrO34fyIuSlKmlu9unyxlTjkubr5x4F9t2
aw4CzOVBg2IEFFzYEiOApRJ4IMYpXxtqaqxc29NKYDvyLIOiIFB5sA2zhlBcYH3LhbNCIQBHoLIt
PqVvlDER5CEzvHrKr7KgqyxTHz65aELuD6ujcDRUiVTLZ9Jr0cV2RWmuSZELJv1ucCDXxgmfFzI1
XtM7V2htkeSw2eb8lrc+PoFiVPBP3mKJpMn6A+HAJl56AMxyuRQp22xcj2dsJYLwfIunGNONv5gV
5CN1asDWiICTSPnVImbon6iOpzeoLxrruONpbYoHui+F8BDdgBeEOzZolIxlehCDDa6sDiUfnnjR
nAszGb7H+z7OuFq0kqeCf4csY15K6UUuJD3UOSn3j/pZ06ctsbh+fxlXlloeM/xIBztFlg01RKQl
0GwrLWVxT9DhtKr34y80P4Gog3tGv1VV3nj/CHWyHyRD8wVKFfnrWjYEd3ON/sgMoKTTgNvS1Uji
sBlpBMJJptGU1iERxwKfbFaNAfo5O998AdLWiztd8bv7e5/+8DSca+r3ZhZQtF02//F+TnOdYxMD
NaM2HP2BW7MLpAjr6fc/ebB1MvjPEXXQzkHuEWH/aK/Joq0txeSii2U7Nyt+3JS//TL0H3pKzzUK
0oijvyr09wr4T0Wj5WBj1r8ha04ILcppSakQRv3iwJqJ+fVPUj4AuWqxj/+w66a2zQVgq9m+1nBJ
Kvmf2MH9FZhO9IioYNX2pY8Nis70K/v5YlUJQ2v5l+6ozZQIMSHwCY11Kjiqdrv61aTzlb0wGlC2
COO0+/T3TZBd4IjwiEvFnk/eoWggM0NkgVGFiUppRwx4grj0rZcygaM8+SiZYBhTD2mYWALynKr4
mWKeFYpUaHMML35zk829pR0NdPTt1zP/rNwVwzXH3hlNCxxq59KrnddH1RgXvyDamgtHd3dJClku
svKNnDA69oT3TRDlrw637BI9uFx8HcE8Rl3oXyJoMR0egVo8X52SOlvs4TQTZsnteAmbBU8pUK3R
wwdQZ174LuH4nL6ojv8pSBN/MyMDe1APba0oCgSs9CvOkDhlGkvIkXkZg6e/ffw9OWmMxRXkWDJl
F7C+z/LCCfdMpEeBEYSWivxW7nM1NbiqcAVsR0PPfWk2DGTjaKhIvk0/Lk9K4Eu96u9MM+vTF5Lu
uT5hevCrVsvgvlWLwd1228Oe3p/4a5HM75pt7o2NQon5p40Op4PYwN/X6TOlCdIm9aPzzUdyfSEv
DRiTqwHCk4UYFlWw0XoHGahJyCJzwFacBrtVQnwdCP91l6PnFZML7eRjw6izyhM57IhNBw5Gy/gp
uPct+Stq000eFc9QUsHlb9MaxLbiKZNGLoHUlmZtRoMuZxIBPmtO+yYtZQLjRl7ROtA+2XZJzafI
wJj7HYez5G2ZlRkY/dol8sVDRab/qAsq4fTYipgeXUrLt6cEbhl6iYaH8OUD6olejTCYz7hr6UR8
VOpAIHCSzKrZTrEsPBxpyyKLF+IerCntBQW44RatUBuXI+7k8xwtRvRxBzt+4mDbvsgCFgmtpbb/
Z3doi2tGlxRmPVpRzEScoSv/LRL6XClwRhbi6FQ84bXELqFjQbg2J5juEO6VljL4A0l9WGRYx3i0
e4Jlo6z0ZwlXJVyauj3jtnVnGNnxi9U7X2NQhZ7Ls6Hzp2UixhMcTfH39XnOweDatO1Q9xRWyJNh
3LXpRK6tBnDEt68M0FFXH35eFx4wbukosgbqGEkSNiQieOJCcb3Zd4K7rTrWrDFb8LtcMH/Vtyk0
2uz24J9b+nyqb3uyFy4P2axXyd/4OoIpQt34B0ThCRJ4yjFjX5/O7+xONzvMLPRcM77M+SOO996M
OCEBNJ9X5DFEMpS0LmJE0sGuhkXSNUmrF0BwoiXrerIcPcMGSW3dP+KsTubAk3eHnKDRnyGKjN5X
Axcg9RmW4gv7ThlmZX7bFDdxz7Yys5oSPprg/yQ12FPKepDZ029AIL2boO+jHNP3lZtpzS83+4Og
k380g29wuezWwF7aEJDI7WQbRfwQhSSZc1DHTholsyWMMDX40IrYqOcp0denhEU+Xab/7tAFCmdV
ngOIVFpE2YbCvDJBCLTrhFJsPbVMGY9LmMd8+nc3r/KGVjpCiCRaTnUkNeejGmGHfoYS5f1mIuhz
tu1xnxE7pEU3zMEsT6WQslhy2CJuxrlryQeMwL2LmRXLL0DR7wUapHNwivImhmj3I3lPRNwiNCff
WaOvWHdM6rvL0HoEDZEKI3NVCr7sb5OBz3Q/qjrum/1nUnBY3cRSGBbbew+O+x0PBJUQkf58yC7Q
dLqc6EY+Co6Ev+Lkt/oh0Jh6W+gTn00DQgT/xZrfTAeeVADEeRSdHbgyZM7RieUrvzIGGOZX1BI1
aHKshTcM0Tw6nd+MFH7HPV0yn/itJeWTxN4yMMlmJ6jpwbpG0j0qAiHLwrZpkXLsMIsIDCmi0pfK
xRBj8qhNXExcvooc2S9fUKJ112yyCGKNHctAOQ/C3rOOg4ZCFqOMBhpQJkjqu/wMENPKWpUwQAUm
Dbgr7iXXTpuUoQtkASbjvcUH0q87NAGTcVFlMS+ZUkcEPd4nfXm8bG9+3fy0MKERcb/RV8/NKpWU
VH3bvb7mXThP2xn0p4KUjfe5l5NtkDA//LcDtAGCfS4tkd+sCMsdNm+MC58rocfsDPkld5/h2Qq9
yyHYztP5+12YTsmFYzKXi1UkORbbHj3OiWkfRgu4R5mogYDgHG+ieBULpeyUCBzVJdXGGP6kSv1C
BZEprsZU2kZ+YjHzvn7NBk6t/CBONGjxTUUaItvreyhl0aPL9ImdkD3qnOIikGDN3J6A5brlcQWx
wlK+4BvghtYbCp92flkIax1n45leOkjhFLoFvAVlzC25RSvPVBfNWJ5Bx90vuj+Syr/jXQ5L08O2
TzitXqlfWOQxt2HCyE3VA8Sa4hZ4FT8zqOW3B1lmekjLxD0p2Eamq4c5hHW3GscD8uaBtV5oD5Qy
rS2SBwbG7y/Dto8CrOgrmhu2sOvvG/BzahehHd8lK2osIzTKUbjlRp4NS1pSxLk+dqPEp8hwzZyt
WYCTO9ODEgVp7tSnxLsPdQjii6uQ1S9MYG7n8+5eOjezzKHwhRZ80vrkWVdjugqg07p8L6Qh+6n4
BDinEwYaWA8du0RcOqnjQrTlj05sH+Oa+uptU/vugoy+QIyfHWncDnNQhJbKP8VPOuVjJSTMe+81
bH5SFLrYcOar6aJIqDJJTzDQpK6fpXv8aYyuJEeN8xXnLQxaLMyPAin1ewpzdpIzkhEsIJY17Pyb
SuPSgpnzhLW/acj1RdYHUdQvvpUjWGoCpAuNIzd2meNBcwfPzf5xiuNR5Wvgo1asX4c0hhrcB4LH
EO7kSNEzMG2n2EahFbYkHADPHY8WNvfBGplVDX0LMu36DHJ4RWnoYXG+5k1J6ANnH/aUqwj0BFNV
SX/PBaF5VbZDfrn61lSM2ZAwV8PED0UKKE8VZVLwiDLowT8b/EAfzY+OcAsRVWBlkWnzYWqqCo92
UTS+Amst0+2JaZERoH+oiH8U+sR6I+CzhtBAiFvdlDJmUs/jgBDl1h+Lg/GDr6bmdwBoAYo+5n5J
1pwe3bfBs0PmEAeqpqeMCWFTWjp6h8RPOTlryBVQfNI54CoK3H/NqV5K3TljZGxizoKi0SsM4l3E
ZVbKdxL2H5cAY0e1gwTQia6f2sUru36QuQ8jkMsvqaNSkQ4vDRv9/Ml7AbSCeIolJ2/+fqbdZjLx
jyFE8qgfE+ZakUs4A6biI7iDArm17iVBVkyGY4/PzHVS88FcJ7/5kiYH1WtnwUsF8Cp5dlCp3qkt
3mIRhHoahIuEUoxOqBzQFCq0nFTVTD/6iwHMYvltl9LZIKdi+Z0Z5lFOKuR2UelQ+cjpKpv7Owv/
7wNlbt1IB6Hzubpsw9N5oNcd72WfcStQQJzZ6mK9on6BbdPxm1Yq8xm0+h7hBMvg34/WSgzLxE0B
SulH90hOioW9AVZEggofVHyDhLuX6S9OqeKrPNJYtBkrud8yd7fNC86eTYUsR1loW4YtphV5RpZF
mNZGinfdkgUgUvXLtpf+LO7Hw3FXA9v9uIdrkOiFWFezPR7MKGIHBpco5ODokFLJJAzLaYgd2883
zpKR3pkaU1yZGbtS/+zbV4a0bvvm9iXHwNi4N1f5EnjEu28OpYDQrJ5WcS1wnAdHTUZOawD7wqsZ
wDFQELIREderc4qQtQq1xsOlPgCQ+8MpzNCvXNzr64r0OQBrYE8DwtQ39+Ws1HMnA1v++kAPq8HG
75IFW7S0qM/tcQ3b1LjBcGItUeVm6bOF/paHE0mDTJtDP7G9M1FomAK9OJYDc10sJatpzIrJl9Y/
jsD+FaRRi17Ootq0n96pZ52PPZzVss7c2XHo1btc0OvcdO6jJDPYKpvBSKeH87FKh9gYKTSLJ6Qf
dyu9ETjRs9sOaNss6hn5Fw2hAqucDOp3wfIxZhUf56hTcOqQossJ13mVYXAVKdqFjKp/K41lStjN
pWvGDLW26YrGGwSH/9Lldc1W6pQ3J9SZquU/6qrQcmrOjnupeAeSvQN4AbAgcwINMvZXkeIn4qc3
Co5kLvJJJ4JphrLy37Kc+pZSq9lQNsHVEFtl8zDNV/gqVVA4NCfCEkOdyW5Etg4gDvbYcsjZeZSR
Z00BhCw7Ih3LI6tMUpLuAydCC1DmdD7QR9OL2W697T7lU+Qw2myQuWaZEV/3Qy11gRw7oUtUlDxA
o56GlB12iY5H4Yrs2rux9UJ7TDObSbjleTDNRuev/Trt9OBkhgE4Sn9fBsmaGBJtKIqEsagX/PlJ
qFsY2JzticWVaHTZQdsU3Y1V9aLZRQcRDHNIfQ13dClHMZE8ukTmsPwBc5wurX18mE3Sf1z4kehl
9rjPVAb4od+lb+wfC/AZOSnmasG0TqYZ9WBc3bUv3REURGYtbOqozSaBoCguDqqbAcc5sfafte3H
XbeMdXrYgsNHGIQ1m58zqM+WOYYDl+x11abh28oZebtJy/cP+h6D1zAktl3hrCaRIyVp/ElG664+
dQQqoSsAuvk4HDHk/KJSWmpxozHrROs9hB1u7xV2MzkULY2kPxLC1PUgby14nYta7IIZ1fEkNvAE
2+14rt6ZjdIcXBca4qWc1A09LSIMCAVJjUA/Y45fAHmBJjngFPHC67EERWktbvaWifm0qAE5GEfS
m3bnjL7GAxJA5O/20X5S/Vwj/0sUv+P660MdBSWT9UXAYEev2+8Puq84hbD6k9Z/s80EfOGKVeme
6lX687MS9ITMEbtG2cgHEJf10P9OM3qCiMCzBaKGNBoQ19bfhcFckemQbkT3vEEnLqk4K6ZQHT4D
hCZO+y6aofyrgnn2DlvM/1idZI3H9sf8vTvxrMLHTpChtllisXFhj9sJrmJZlKHfiDB9DGRvTfEx
ikuBnsGsqxybwdcjsuGPVGMmNDpiPAPVqtBjfv/vEzT4wwxO1Rljou2g/X+kLIliJVrdeRtgrWvb
sioB73bOz7AH3MH1qZnQxn6+zLSFBcI17GPx1ULJ8wkLkFy1Iaft9KhqzSWj196mBqzRc74nZsSh
LynKXKP6DBywW8Rbm/cgP/BJ/40jIvejIQjI23UDR5liGY3nT/hE+3Wnzr2go8WFcOtFaRzcm8P7
34H/Eq1tsZBOLzZc8qYBmFB5yYhJ72YEBtNUlrVmkB+xsNiDE7gYI2MTQNjoyGTJmM8yOGIXoXYQ
scriB8c3c1aBoMze949Z23Y74x0gNJvP7g0S9b4ipCbqoTCBa+eqleIYqSZEFAj+kleGgy1oNsdb
l2fkiyXsNHqFTAjVx9JaPfWyC6OuyexktoLgLsGN7CpX6itUWKTx/ezUjKzrPcUSxKOV+eUSqjfg
OIz3SDqT+Vk7Rn+9ahLPoCFCpaWGYx+Ao6hAL8S0mTfqDpKeI0bD7QwZ2+Zppd+wnBKh6DtI6GAO
zCiPu+rKbDFzSfyeScahdSxgE0qkhUgQzzXqA72wQXf26uUB+RFabhVqLnxBN2U+xLAXxjqkrBlv
L3yHcWICzKfsnXhPzqSwkTbmriKJoPNmatMJqFmHuCKpzU2RSShFQznmJyOPFhYck4UzBKL5xzb7
lJQ+ZcXK4BPAzkP5SqzfUJ1yz4qCUp/lIcVL3J7J3DRoTKYK2e4ARIPPe3i8pDDq7SpTQxQlTaKm
mtENITv6kaL0l9A7njykV5LMo1nUVnjzouXg1AApkwDv8uOx173a2yeQo1y0zSzc9+tXfh7Ifnua
nCSvDNr6/PJ5tViBaf6YjrWW4dtkdlxFKwvhPY5H+tgY6VxCvqrURaoGXzDklquNEZ34M2nl5xnX
crE5JWDkmSUnwgky7yrXNzX7KoPkFowL6vf15xbtW12z/DpdHVNyhLNgswFDMidKsJawadAFBSEz
XpZvYBot8ttpgLS7AtyZLB/+4qZb/bWwR4ivG68lV6Ful5nUGCXJg5yAxxhY3OAwSY0yGn9ut81C
aiOTwzGTol6ipu4REUO934OrjRq7oEeEfDwPSOmq1AOKzFw7vSo4YV9OA1PUu/Jpnk7yLvaRpP9O
nKDeaH/LMRQUuVihoZPLChkAAPAO9EkSwm8TgCx2/hF+jBMsVjRldd8DwXGuIkRGXjYGN7T0XABb
ugGWly/OqQxu2Lvj7qiT1TiaOJbH+1sKB58KJtT8bMXaYR9ZORM4CGEP/PwaoEohRuEgtyPKXAqk
d9HmTgMAoKJd03f8xLhK0JH11zqIeSSbXsN7e7LCys+COgzuiekQQ/kMtBvq+evO3Ak8vOBhLRMJ
Ugw0uBNRZ2t/ZDvIIs/nnsVtgiTpdeRjXBZnReJ1u0Fq1jrFeGkLpSX8ZrBNffy8d4ZRvlW1n/n5
cN1mBMGYLHZms/7EqCOdKqUIkGQz8EHcjnsGxVTz5LFVBiWoOJMG2TWUsl5DisCRJqbUsAN+Dll/
yvqG9aZu1S/Wij5CTkAAeW0umswPWf1DMQRbwG9YC2ZToBL6HjsobOdwmmrEkBxbAcOXa2YbNa7/
j+5J51nZA1aOJtO5VSL4sS8BdYQpYep9XUzK4PB4ZAaYV7Q49nwKKpafm4IEl/6MKAel+x8LSWsD
PqzX627fXFi5lU8DexGTMHOBz1eBZ2D3yN+tOy9wjLXZI1eNITp0NCCyDCEWX4t88BstGnlSy7QR
Rtu30FSXKNkUqSXIpRWx2KaDKUOC76X1YKqfBEfDRhzac8iL5bPOBAbwDXxcxlLZ2zuIQN0ta5EI
oMZGiTucLQhLIj34ZrYbTeq3opfSjHgSSAtEjcFMLc/oJLiUZ7yFqvIn4qeHaCN7ec/dSrgiSeoT
WznQtDn3gcavH/eRYY96Bttnz8HQ5AsyXIkrKMftKSTaGCPdlc4Rt0lzZTrPddlQQELotrBNFDRA
XwqEQzqE/0nY17NnVyh/a2GzkgDXyhaONeRovbrQ8rKpi7wUcUHV5BY43unIRVlQ33QwBr6WuPsP
3Gx8XRjg1ksuYTy/ITyOpjSF2Kgg2chEyadrLrova18Yzjfyx6lUodzpRs20gnTvt2u2F2gdnADo
OkUp1hR/rPcPyMbHYocuXp5piFHa+FTLy/OBM/AAs6MEZGrPfEAc53nbQNngNHhFJhhZasXA/wna
1AE0xzxhf8GLa3jEIYCMrJ5Mgfmr7WhQiDCUQ0Omuk/dL6kkLaZVIPOfob8Ivy1zq3j65+qqTK12
Pve+0Yp+zO+CktkReJdgD3fzyC5H7XAjxFLP4avEOOgg1sLJDbLc8Y8i3em/1nlBgh/IHnVa+76n
vpmorW6bVHf5kGgE9ytCgMxnUKhSk0rV5BI2ThM5GlEEfxwMKHcC+eqeh6jW1HDd7Ao37OmcuLw4
mZTfUL0T7HkIzENTOwo5caXUuLN8FTfpeo2MqqB9/ZXOIF0lvMOVoUfUt9PwNxGBIMQaFrh6jXKb
HvbOAcj5e/JUWPI2wmbfzsKC+7WrvM1jhOz4hT/5B0mZx1MCFegQfLJcEUXwwvPx6rwnciA6b3pm
kCQHb7UF+TTuiKVJ0fvswWW+dJd07oVhULoQg3eGqnI+gJfOTMI4USYvJeII4s3so+E6US6Hf7Pm
AUM4i2EMqH27Se4BIC5yWlMUKy+t5NV3t11B2UGbgpM7bmszvcH5vROuJz2YPpkUz6E0Vx0eVv5z
v2SHtDyyt7ES6rnblIdifKmUV4uQUKb0aYDvKET4lSgRpo5f/HTksX10vt68v+odR2x+5XpdKyjV
dYwBmjqx2intSOx7TRzY7zzWt1DGbpF7K4dWiiPSrmnTH8PJ7rfhEQyljgICm0m1mM9YoDOmRs7V
z1LRC09oGBRRPNkXnwQfOh/wJAoibzxw2ZjbANCe5C8B3N4/A8VRkDGtTd4aqr/riaCF/f7Q340l
EIxxvhbZqW488qis9r+ZPC5iQoL+H1IqHBe8re/w4ktJWA+3UBnwwdHJFOu0DaXkhjHtHZlS07un
2bzugzaw0i08b9mIUo5mu6hVhr0myk+EU6ouoYanwzH9pPzb5SBQb4BePXtxahcahZxOSItuWFsn
1n+/3C8Oiq5JxcuwxD7u28e3pAmXq3ZIAyh7Hly+hTTv6JGZcOZJpkMp3kITOuhjq8X+ye6c9N/Y
whSYC02hcJ/iEUyXJ5AOAVLNsHfnX7sspUSQh1nczsUjx+ezPoXn+2CG0Xif1RWw8pitRKpcN21p
wIST5DcBYtrZZJrE4AzEJf0bgGlgLiyVoFRUuxd/ijTzWb8KOUtnWpTOcah/zEZwEcCGCxB7pkwj
PxII9T3j5ZXFtLg1Odpml3qUfpHn/mp+wZTxuQUbNQLRP9yj0oPSQblH6IPWb2AtIHNt31BWiqDU
xcz97HkAktVO26JvONo8EgQ62r0ymD/lhCjer3/9HurfvYcT9Lzvn9foXINwUjsoo0FPBKlKSZFT
uagshjZUUglwc3HSrwJcfpiMnqHVcRqb2ddjSZDrzQTJpmpSHcpzvxTB+L3paivjipJjKwerv0qz
Un8bCmRfM0+OEpPg51x1GSlAzq3hbq4s06rE/bR3FHXKZZqamHE06PqdZJFFgvQbZpEedTcYm7xJ
BYQ50l0MIdz+qi9hjW+304Hvt28Bcjg909XU+Fz5539MyWEdwU0Iy6joRYllUbUrrIBD3RhYnm5C
G/kUqUSImF804i4v9JH6AEGVCo1TZ2F0L5rno0KdKBQaETyLcw8uCISX1roB0aERTEGmAQTFWERO
+DdL+kyx7AjuABv95b+cGkoLiiDR77pN3WIFrxWQOHgtPJeAlPY2PfpycP+t+gKNxxbEPPHerK6h
OaFP81+2sKsDgoVxcCE1fOQjojc6aCesnaPpIkJwUhimQ/yacXkVkLfLhcIvbJrIWVa8q6aBPScE
ocpFiQCO5ItZPe5vtOvC+ePtfZWYSuOslTTJUM0rtUMgpgCoZbb8ciyrspEdKYURc1lnwLyFun6d
powwOGItUeUcDyzPOG56PjV9RSgToWSzAlN2RyBT/S8BdqUzlZedrDv5I83Wda/XPHaUIqAshQrQ
8jn6L1uQC5V2umAmF7IJGJnTDrNfvPM1l3PSigO05M+l+4xsfAJMdwXIrNzIDv4cgl1xw0hphtmB
lnZIEQ7UveKbwWJzLl4UsVmsU0X1mkhz7p+ggFrw5rqR5APv16soJwCXzqK8Rg8VpzL8lUT56n4m
vBqQzy6XkY+g2aIx4mMRLp6VwUdA3UB+XgizvuF5fw2GIE3PLNp2+VnafPj7vm0xdi1mrOY10Zey
430K5s5b+DR4Ef4Wlc8YeO8B0XQXFEwqLpOXf/f47KhX6WKn+DGzfsgmjhJTBTgbT9sv1CDNk6Uo
XKBy17VQV+C7sh8UzuHpMJKIaysNu4YqTLgswhR9NJCXqcTsQcno9F8nNstbF08VOLRNClPYuZt2
av/u84O0Uva4JeHyQ8O7xCdRU5prDcIefhd8EResbLlk4qeSdn3diUpTyoBem1GTwQm7fqQw4tbl
/UKMUqzBdaaHtonjKUyNvhD/Z62L34fbP71I+HJH/yxklFN7isO1K4h/BKRfI11XVkbdO8+qItTb
dGl2tQhQbhpanEsK/0rDownq2N1dgZUyyxXOtRukqU6m0jXj+qo//JfgHIxlrBTgAiQvL6VY3YTw
5ATaWY7AK3/HhDQHj5/MEROaztJPR0YlnkioRtEH7TpKSTXleLS9UTU7jAw0bc8Mlb0DTv23MP4N
WzMBN7J/GS2Glp6uzV6hIBIAfpPaWQF6nEg1bDbvjJxZikkJl216idgc+Rpp0+USJ4z+aogrKxSr
xX+LqUW1EmFEHDtdzspfSU9xarFWE5VIuba6PTMxgsrmRg2x9yhrkDNp5YstlG3eu7IlTi3CTw4w
47IcUqUNzaUeWzqHlao2g9xS+QwdOGBdSYQ1s+I1n+VweUzPj5Gb+O7RaZtGHKYeHr3QCuuo9exJ
va1XmgR4BrMn/yqKFrPdzMDaXAYZuBjvy0ebq/v+ITrGDopgRnFNdFOMlJ1J/Dil/bvCMWJ5vrPa
0h5MGp+HJ8FRV4iveed1tOTwiG0zpx2aUL938Y5IvqFmbV8mkzMbOjceFk+2WrhcoTVC6srKmBde
MVYZhJQz7aK7r/M4DxWm+vtzbgJVkyxFYaC/g2oaWzJsMOMojVEs9eUuaxGHHKQXa/aGeUTp/5R+
4YYlgfbrsb2epLs7TNFYvzXcHkGVbQJzn6LrRo0MF1WHsxRKvQrzzX/GRO7+LWof3qZEYth8TRb8
pSM6rMfw8wuqP+cM7fUhAKW9QivTawEFiA8qqmZ07GhUNki32MHm+HiaDPrUmAUSslRUk8Hv+WZ4
Q/EQVn34UkOFMCtNm0Z3g239AniytJHZpgCJee/94GowJVKxl/bk3QM7ca5JnDNVj3VOAVS3f9V/
gf29LgHCWkSITZXrQymce0xShXNQZI0ga00dqPSm7nUl+E4lFstPa6ERmCuXqQPMNRijIbJblTRG
NHkeEugxo/i+ZQi0AU/mD7KInRZlsL6fXAh2xGNquZQYlp1vvoB3dFleDOOry/f9D6KIN8rPfgPS
p0982h3xFzXiQroxi66sVqIrm5/kV6LAXvU+HrjvXuOUPsc+dxMQikRVFQ/Uod+JbiKXZ6JDAHB6
fAXNkpar+HDXG3zs2wqz7Bh4pte2F5NiS7johM0NRboZOJkUEeV/w/PUJbC4smQfNmbF8uxlZqC9
ONs6LW1nHhMZt6yq/eji3rCO88QA8HSLJeQHw/14XNd1+dbAE98/mCWdu1jQUzuAeBYv17VFuZo2
VQpEyJUCqisj3Hq6OQWE8bVwev+QxW44wcPT4egGzbsjo6+IRi3ouR9sgwvlLeuxcgebVt0GMpG8
T2ke+nBrrKlCJbxjOjvtURwrWpJfhbhkZ35GNogPudCHDsZW2xBTOev2YgrrvnsKx2uvI1vUHDtN
AmiorHo5JYk597oelVULDNcSpT0cpWBB+GRbiWKF1LhkhnhchsrBhQnm46rMwYrgvJtWgi6A5H/Q
ogp+xmINkRwrTjem3Y5PzZbUQWwVACiYJ+fOpPK5+VNYXA5nLueoZrMNgHYnmVIkE7tXeAvx+5Md
cUp+xeecF8zc/+vxM0EggE8RUNGttXyJh3OyK/ZKYNRflPMcaoiyg5O9PxrdVivtXtR4FAiJ0+hz
r3eryOacCKaVDQPHuVS3lSnshPPWMnU4Nkv7M90Eh1WHjhHxtmNYWAZC9hZ53iPPhDOpmcp1fyLa
VMzaGl6yoynikaVQEulDZ+ap/+7Bbqx6PrXLqqXdgMMsHLVU95eXO+XRUMgnDnmjeW3WA1kRU6it
Kg32nuQqHw4HXtSGTfAaaZwdksXRry3/FSCX/XDbSr2PRYLkGSrq75R30jXfUzVUwRLhRSvDtM7v
n9R/GNsnUbFxLJp85EroYE5mMrPYUi3oa8gxH8f92P2QD9MzbPQU+fOzaVj/E6QICVEyK5VR3Qol
TPVx8gf1aAlV1n6T39bPbnwP/zzlw2hY5BO2zxMp6Lr2WKzBGQsX0PKCbEY76AbhFJNwokyQ28ou
rBYXF0phNuKQGpZMQjmCOP2PbK+EwEgTV7BmPWUD+o3rPjc56u14VCkcWH9DuZ1BaQ7Q80FoLLLm
hHO7T33uwIqCv+hNJuY1He3GMk9Vq9uwhsv60kMRWRejRORmbBJ+pqpwLOPK8qMXewbyii4i2LEZ
FZxriD4BdwVGIc0StsO2YSXs/PvF094o0kE/dYExq2jVZoWM3od5AJcqlZ4V9NgBH5m7g45hdXQq
bQk+2YEjk6Mn1fNjcXjR3k4lfenBXW8bCIWyZDEc8ZEzVjPFcKBl9PuVW6kiXzsoCUTBJ51bMNtl
qU5R6JjyxxhKdSSmoxEYKUCC3ksbtN/yEPRM6Amu/RT2fw2gkBORg93r71lthWGpYikqnOO5UFXk
nLUZKsWeNn3AHeLjSzJG5+eVrf8QhMPkc8eXyOJClE6Kx+W5DOIN/yK5Owbn1wi4QWjkzuY/pNNJ
listQ0QybJbb/yVmfS+9gDxb0bOJogqed37h14kamV99q0rfOW+nk5j8Kth6C9Z+woGl3K8coU+7
0NmricPVMw4iP0m3hK+H+7lol3i2nUG8cyZ+oo71JIU3roGFGaps5HVRN4Si3CmCQeqiWQ4FfQeK
GjPipVkMjHiL2W1E8UzmfYPfGfYu5t9pTJrU1kk4gkL9tfiiHPyzMK16T2dkWTcLPzZoVC3FU/QL
CPVcp4sQFtWVRiVXFivFJn2OBb+oH03BEzYcpUc6bvK0PiQZzbWwGvKrkLcSIUnUtpaszfNyxhY8
T1xH80sfoniS2V64AKZUcXmlyu2s1vkjB5SSGXBnzKXw7q6BMeRrsdNZt9i84UQOFakT1zla3qny
TCJbtPhFELJmiFihgP6na2tmv7PppUHUYrxi5ySP/rIFTKL1q/u1WLn8644yQuDM0TbZaOEbuS+q
kB5bwnUEN49s/niuJ1r82lbNEISJjt1ot6UgMoIcNwoOcHm/lUj4KfrmOAnccFJwdqbge4BPbdxf
xe8i69oO2ASdGVvcbcmphWkLuTw4P2Io/U85jb3nPYEGWtvPoqZtahtRz+5rZyQg6QBb0fCqR/eX
HOOqcDhOes7xQ7g8pWqSZbDzepO0m8VaECoWG9FtSSXuPLqgJCsO8jS6tCg2cfzEek9UBSeX+k4E
QsTzBF+/eT+Za1W5g7UmHZ7HUM9cHfU41Pq8B53RNd7TidRTwwSCKMn3M+AGClCALcHuhjNCfxBz
XEwSlmWAKX1zyKx4vEweT7CfXPluBUup3eZGAb5UNkeAn+PJg0QeEWkW6Oa5WhF3u286nWYZyYZl
qFmIepxbuF2r7ql3IKjRd9Njd47wtc6hVGkM7cG8l8JhEJyrbusPTNFI8ZmJT/gocTa2sbdL0Reg
077iYpvsulk4Jei823Ep0w2T3kU4tuzhqDGV6Huq0xWNlxUzWTmjsc5xIw48nIbWp5ySkLV16hQn
HZL/SLOTcpRK3xSp3OLJxdODv0+0fkCFRn8yxfSAO4msEQDxdHPzKejbhML8QlQPxfl8dHk3f7wP
VMc/sjBiRZAN9J+ke/QJG4eDBe4gCNRKM+FeJDSkWzajYVgeHoDceuyzgskgAhQTX5ojuXJXOKB5
dhX9ITc1jfb3LWp+viGkIAbcPOsY5uDxSG9zF0lWi9t07ITCSHjHyZS1BaR5S9B/GyEKR4eakYsV
yGcuy4XKTNjTSUR3yT/cwWjNllgwAnQOslHBs/o6mGG+Y8nqb59+KJBvHGew2jN38h/5M4qiQQxy
Jm2yNB882a0sxwuKX7JhJEYi0K4pGovJ52UGSZVBeFDDKRSvu/K6pl6Q60mLTCelqDHvzgMQxJJX
NOLDVcXq93Na5jyKnusJVv40JE7NvO2E+31s3iTC1m302rAALM59kopE5rd5/GwUaaShtNXcDo4B
ed2Kr4kaoXqCXJo3Cn4EdKr3rd658jqgxXKQBKlVQh0PQYR9aEbK5kG/gXGPbTKIpcLFbjgMEtlr
n0QLLgueGi9LsjJ/kCBxv1wLBdnDuC5tc77tjgShP3ng6E4gC8rX0MJIwpv5r6HBQfEozr/oaTTU
IDMxT28NSDAkUOuCVCTPyQLk1FvAs5nJYjWaXCWkrP+CUCGnFOZUt6O6yA/MQAaUzYfau+8gfcFh
IXkS9t2tJIajQz+47P4OBse0NE5oTYqzR1DJtWs5/xSoIfI3D5g1wV0NAoAora2ckVus4sV8fWqO
+vwELCo0g2p/aacM/feJJ6CH0RbUsVQENnmiB4CJ0JM0oZIa6V2obeAq/Yx9/qMYmMzIlImk6YhZ
uo/D3AhxBm8cuAW0ZgGBG14vunCWhCtjcpNaWmdv/k7Au0KRH53iZZeQEsup6zITj79o93iwhkfL
4+OzjKgEXAWI8FyeyuXts0+PxSbK4+vpCG9oihWt8USuFkKYyXHeO9gp82+og+hrJy84ZswilJ9e
Jvn3xjsDjR1RGSVOtZadJVKm01ySnwNwIxd+z3VyAz05GNSKeNCUIHThQd1wyNPBsKPbR5d8aR6v
oC+W2LrJ1kszLjeryuB198QLHwC6TjjnyvpBHM02UaTe6nS7xxL5OmpFFHM0cd7uEHczGjT+SFKS
3JBWzhwCXD1ftcsSgTGMnX50tGHHfibYyrFsa44AThFlOMHRk5rgTBF30knbI0DVsluAI5eqn7hy
RjCoMT2VqLK7kqp981TAwCtMskvuV8ll5R4oCSj6PIjaQaIL9KwF+P/COV8Hgy0J7ntgcXtej75n
G2Zk6u192AVRFm2tLEkAhU7Pr7d4sOELZ5ev5PMosdVT6bckdpA6HqAEVLEiFbwg/m6NivqiQZcb
qyc+vcaDjffPlVSSqLfLnMpuRt9gMDbIR1tbDX8RHQoWplT+R5n25JBceDXiEFu7gSBvWIeHX+fp
uwZQ7Rrnmm31mmZ9h/rUsyEySDwy9xo5z1wEPU6BVRfNCn0QFrj/lgFEGxWk9MuN8EupcqPtxWMS
76MPQzq9COj02eV+Hb74zx3Nm4JmTvJ9m+yolJavFDgc0A0RXlu5ARz+1Nn8Ath7PK2htEEnLmgG
+5NfvXW4iNBhXmCZ75tJN820LUkc8pCWOonWDF3qlswIze441/tG1dnKxDepAVbQ0l1qdW+m/ZYj
SQvPb0uZDfVNj+tjtsP1AsVxgxndf8SiAMMCVP9DND1qIUazUZrH+FFRwre3yZEbAywFV4+6c/dN
SzkyGuTV6TErwJOWpzbCAPAMa7QQ4QTq8VuronBUqk0isOvqLjwRSWQ2eSD1de6qofdXQ2bxMnIA
q+BUgFZ8ejbhtP3FGHlzMZ2E7NPVvzG9KvI3EsnSK0rinM32vimQmAyTURsUNGeXZnuj0PEKm273
ahto3RQ523zAlvUH8lnANpTJJJz07bu2zAoHOfCl/7LtxiiLdUADfXDWxk5StjFN42X9KnAx5avk
JExRQAS60j/werVcRVOcQ1B9U4yLaZitHDkPM5+c0go73jYVH7xG3R1FkQSjr7+4EIOYbODdiLBQ
L6qZEtLLMzT8bfrP9BPQa+wlsJ2W+QtxPEfcLbmmYUwfkPhzEsadjQVjm2XNwWVqGjkyBR4W/hev
OQUFum+o/sBQJoRmoxX6pbs96H7bBS71RudO3q0DRkYIDqnxYXTTls7VeVz3y2wi5j8Bnog0TTyo
sSk6/9GuvxoyYTaQK5UpHVtx9c14X4Xo9KDQBqhAonse1WQsZFCqaEFA3SQQoDsvbiJAx4rUmk3l
HYyvsbRI2gmEmZKlWRlsKdvN3rDpSDm8omphmFx0NrXDrvlgkBAG1bV+LCMqPZFP0EpFZjvolX/h
8/XfPpWIPMBKLKm5XdRPG+sFKLizZ7mfUdJFKIO5NIsLHH9zPzxZJi0/sWTJ1ClabuRSBq9LA00y
EBY3qzPZBSFMPk+9g/gPcBjN+I1hAx570865AFnkHoiEstdr2nrU6NvAh9UQDcvD61cjyCM260ea
BIKfDq5mZOq7XgN92PsjxMG+N9/VdJ6W0iTixtZv5Wb5ckdrMNj000UMkODuJEJV/gSZ5kbUwTTI
/7v57WaZUNkczbGkrFZ8yRF0P4493gUBHqSPKzq+n2leNtESmfI+PAK74jpgkcrFQLMM7rnvJMiQ
dl0OFxc1xIPv28GkoZVoiexL4hQFBfPc20FjcXLqTBW8lrmOLvifbMbjqz8P6SlWDvdBV3UopkEd
4yv16JttDjX8fBHQhFLl9pnIaSQwVSF0Vn0eo6cSO5vj6/GO6LS/+vVVcImT6DB8aakLTzjlf0tS
QIqkHM/NXC64jH6erzzoxuj55grd28xEMJXigFQ38oQsZYgRx1nyL+QzKZBgF3LFoMuup2rYBVSd
QNFtuXceT6bI1peOUbQYD2V6hCGiuMKlT9DNiMYN2rGqp3sQT5w1x5nLBeKNhoSayx0nXf9V6+uE
ltEUOsCH0CBlqd3weUuHyBzPiVu/ceQTOzBLOa82Zb2ZaQgIPHvp6BKTfv4tE+L1u+lksd2Mck3A
WKdKd7lD6oJwRgAZyyfN2sB9a+Jl/x1NdnLFS7KTBTPmOYAte7qnJpQlGKJCG6ENfhs2x2D8LY5P
uEwGt1hpui71uPJhf9g+hiu5ClzC2PrbDYhrOFUMoZCkt5w3Rps8eZL9cLgyNEpjX+gHSB3bC/fT
Vtfg8UebhscWBiRvJZlnC9bxWhl69k1lrSGwZOWGUjj5xbyZDqzsTIvjFZZ6raE9Bgq9PL8mxAl4
CUcEpMu7fTq0BtcXp24q598747yWQRhe9Iy4Sxj+tQQuVYHcmhPBT9rlOQS6ze3z3foj/ztYZU7X
UF10AZZNKByRBgj7XecHUg1ZNFrD5Y0HbsF1pELC2HEuv2G6KavCo4PWVM0g3GU+khivRJKSqLtz
krocEzcO6l95jOe2jtF2z7IuvZ8rZwPZlRcvXckntqBGWuuln05fEB0CXFmC0/8YWPWU3V0HnFXu
twWcMeHBdv7Fh0U2mFgaDeplVFiHLbLJdxginArqnfIZLc0YznWvOf6HXb3djA1rDlekQZ5c+wij
ueG3rYi/HsunCtpUyS04SWUV6SiqpHzK3GH7ePXdIESsPW6qstbTx2KIydAoMcv81JHZiK9UbwO/
IDReuiz0jUtaRiVzssJEiLv64albi7jKavTw99FpI5PfHv+ZWyDU+H5fuHruKWZmX3cxhSO8F64h
mVv97CLfhpQlXXh15+Za/pvX4WXPWG7UOfOzth9RmlGN5a34vW9wprc66l4TKfldJWU2TwDNM5Vh
L6VNXfOAZLu4Z90d3F9C3++xs7nWW06wgE7jEuB8HaAsyxl/kNIl1QuuuIrszLEp9z8VfL6VNvBK
3tgeEX1EprIWXU8NDoEosEeQ9kT2kMPw+9dgyA03tWHHyfg1ZyIo9V4oGFaVNdesxEZkYq5ucMuD
zxE2wPRtPZOAqXPeqC23uJTnuuVYyx5VQCwg69ysrrfclx4YdMKQyKEse9bwM9fGUNl5r92whIPV
8sWHu2c6SjU8BhhUyswmkq9lvdb9f9Sk5skHI5CALR1lFrTpugr6ZbHSRwbo6z2nL5X6drhw1ofi
OrnHdZUOAmC0Xmi69EFc3NRx7PR5KZ7MgdrecNV2/L9Wx9hbg/VOm8lWvh1tjx2buiAlsdeCxN4k
Am5SOFiLfJIoFn2KUq3An2IYVSqdBa7QPF0f8wOduwFdKgBrJ5OiSGSqJPa+QWro7fF++l3u8dIJ
hG65Ml/UMEijjIM8hq8A3VYmi8RACSpbWY83dZHTWo3dVEMsHSTRuFyFcImuLSnO5c6ztiz/oXTc
vTD+oIafJToJGxHgCXGhKAqwPM8EYyP9L6gcxOfwuTez0jF/ath+wUGwEXljEeJr7famCCyPTxrR
UUAuHGPCh2wQ1bqT+EvjNqQBiXVXqTu13g0MpOP+qze3FzmtG/OGQF9z6o/YVps1hCyFn7TK+vEr
Puow+5RUwY4J7Te3kVJetHqd3FYiAAlVUIRic86pdFRu2CT0IO7Jq6JZWHIgVHpimxJhxesLmxFy
9nu6IabPNaSowffwHi+ai+IduYyLCe57WHEoXSC57tugX5cDNzvoAM70rWBF54U7vQ1ubtDFZTtz
T7J9WAokRL1stCjZiObqTZDO9qK/WwmKjyLUxg6QoSaFgTMcNhJ4kmpTV2Hd1hPsExKNQr8czIr3
oLKEZFJ7MSNiTflmk/YSf7MyfCXtjcn58cZoJQxoXK2up3WaYY+ODY++1yahVEfqiUK20et/5nUB
tGvnWJuF/hZ/32kp4Vz0KvZZzuQJ6mrVQC4HbkkR0uz7vbtmFKzq7Yxgg3te5w97Tn9HMXPULD4Z
B0meXNS1xHzpWTK+tMdom2Jt0A3BHHhIKDBGlkRsHluX6PYFGJm055IUxFLPmAmzHBk78KkxYCHf
VVNz3TWKPGCwxMlF+MR0xdFcaYeuSv/wH434yd4YjlJIkbWKaSUcxF+6S0dekuq3/yEdX70E8lYF
kVw/R2aq6APOxhF49wwZKIcVhH72ynDdZ0jlfDnhDIgRanRKjQauH5sy7NVx+mKYu6NvOJu0muLS
6IvkA5YyuvYbaOVaAIUFtWusfi8BXzhlfc357YY5pFPBrG18KGUDq3JojhIQsGxohyTj55FVzABo
FO3dqxu3aVjB/o3eOW0WaXRo6/kg4LPuhZ+jahOEYL6rOYm/DzXcS+FHs3w0eY0V5SsFOw+hgGXa
gTcF8hf8B6mvC2vkNIh6VA+GFJlb1Xr/U5Ik4AQcfFaHbNnvP/b5bxbNCuTgMmS3nfrB+cMV3FEi
JBE1jkQ/TRrNUNMyiA18U5WD6GOnJafjZxiYqLnrO650hoX2BcvnWa70Kc3URE9ZJi+FkYRYqJ55
yYtItur4AZZedtJj9ilJMe4Tj1tfXn0MCsREdSNRi39vb7Pg0SJVHEEe2zgPQZjlvTRUJDXUjrlM
TufZwaVSy42cWzAflQN2D3GOX9M/xt7i2IOq1xaFgv/ZK+A5t26tAAoOYgxhnP/CKsHvaeqCfWSE
G2B3pxpeI0DcV0PmSsS0Goz4GlGbiCLgDh2Gd/+GaYI3+BXiNXcCgwCu+R8By3KLUm51WTJCMX7E
vMSbol9rPbrig3YjBkbydyWu003XIk0dmfdYSgqwxAY/PuqNUfJHC8Ev4Q+3CaWsaijoDO8gmZh2
m0T24RTAvSDNjUQgkn/PnKE2zI08y5jnOgKF0jf2ozgwe4fAKNBh4eWfXJdPZoglLl/lUCZ/HdNq
PejiXGRxZextQRmrkH1PvK81DFc5jVNvwYS1YHsyotvPOgr0QxBOfPpKZ+ZOzmSJ4Xi2zfix/mIJ
AtiNlRhgm1sByKfmAhC7YVlzZXXJ49+8cCusInxXWh8clsGECR9SLdPi7SLSxBhlIuhNzkV5B59H
7HF8CkGUPjmK3dFy6/e1J66ykoKT1cdVPjbIzfaxWMkt1BKRIFa8pAG9wcIVr9gQTnJilHkqciYe
V62Hnq3pGIar+eJEHhsJFsIL6MfmW7l6rEWlEYSsFG8bt3W/sFkulV814ZkBWbx8Xy6ngiZk0cfb
KMA45XtFobO29wD++DotdqlAuezeNz3cA20W3nugKLL8DT406SHK6GD8+aJYSfL6h9U0EGp5JRS6
v6Txy1+zgIz7Ck6y6J2mfEFYO/c7FVrhy1uSiSsuoeXeLQ1YsXWRohwbYDlgwv9RZoAfetQEivLj
yujOXPbUdeSk5bUvRu/M5cBXIL/uW8bACN8L/wRF6j1t4oeL2hMrYZfzrXh2grlpLiaggynFXybJ
Z80j/Mkn4oW/RvuiK5soGU/dkAIySYpv3dfNiYVADxbmyRe6wgvHncOrMFdev4cPrnLuiMv6PULx
e+FpWB/7jqXnr3aJWWxTvBzbhM7LbuBu6q5V5ZICSj29Tppie/yeg4NRDmC4rKzSrwC6+EbGAfID
11preOsfiOpTcfmz9beFz8HO/Nz0vZMrLcZ4QTCJ+96qoCIOQvLA10j/+TMXb18sxbcWiKl/A9c0
OW2jY/IR/2WY6GAtOyDGFCzj6QIh+Md2fOXJjJrT1O5l2lPA5I+Bm/rA2JaatLwJd4Xn6lSnBSHL
pm55LAODGZDYMPmpKXmMVb99DdAAOLuaPnMv8mrDKSg9oY0c9bMQrWPhU+Ill+3F1ho7ERIqpbVX
3HOxlJHBkCYc8TBfMhFhi72E2tc+m2/nq+mdVzl/5p+ZnsjP/fUMRj/lQgOtYBJ7sIq5dQ680xoU
aYae1Ib+jwm+Tl91CC5eg+CstmxZDQdq4YlRZzhH3QNcjRpQF1aXau9J53J2fGByIqtnBIz5rucr
daSGtPm7ipnQ2WE9gZl2JHXEB6nybXEl+LJAIWBCxWO7MMlOiAYO1AvEHbE96Dv3vIHM9Fb+GMbk
miqRXk7XCSI8IkVx4ySn6jsfhLAvx1HBB2SjNMsK5lEQhmqLEPYqZ4hlBkUe8nIWbZqpkWCDp8nu
U1Z3eQmi42CT9oRg8xQiOybvMUvNlyFzhvkOafvR0RmUHD0SCW3wyh4NC3dDrSulp2ks0qCx4oCS
25s4uppJaCJIL8d37twXp64ywSS4YNv75+s4yIUweCkrSg8sr5Yh41WncWBQeU0F8WvTPoYZheBp
JnE3LGd3cim2J3M1lP3gaQVVN/NSrQNYCWgfnMnvop1zFnQlRwHFEzGsioq9My1luxIaBjUgkgLx
zv19YLS4+ad6x4Iz0QFOeTkGfVC7JL/Xct7F6TrlmbjjdjQJFSaeiVyaymc7dVphBSqInT6Vdj2w
xVPFApYfw5v+omubU1ifv7IDO5cV9mAa6HAy5PeFRUzk2vk9OnxauT7cnInXcnX/4/r8hvVaRteu
13Uv4t39t8MN6TvzkwQzT3tqHYdOGBPoHsqI4Lu5R92d5wxLvFNE0/GZuE8pT272zWYvikapzoZD
wL3s1ZYCa2+BqQjoi3z8L1OmwnnV7HgzWjngT6r7cgrjDAFvKoEB3mQRB/H8yJQgocZFQpXML3Ms
XfNk0eik6FWwYrfWNWHudVb4hf01aCzYiliq8nB70hsIK48j6Dg0bq6qbYpVuGK3du+c2LG0nk89
VfpUuun10pENP6OkU0lCDMOPwIYwiKXBuG/Lpgqw2S6fgpV7pKt+kWKJH/u0E4Vx5UpMy+c0kb2m
Shq+Bul0HOqEF1mpKn9k9JEePMmG+x+NOgkseLaBEdEInu9EcN8Twx26maUOS56d9aVxYK/rXL1M
C+Lf1DxeeuKdxIZ8cs/xJD9Df5hMhgxRLBSoSfNp41aO8kZ/FFpqvsW8MdSCp3av5RYZc2INOarp
nM+/DNe9EYcgHf7CV6vswOjAJ4/jhdlMglwlhMznmbj48+MZVpGrRzv9amy3Xg0QWSpRovNybt5j
DTjHRv3Jy++iWZxohknhZHlTSqwsBQslGrvFDRRHlZTGjdL5p93RHZCm6lUnIBHGSGTXheF+IC+5
HiOyvITtsC4YF8f0H3ZAmPEQgfsT3GnbHZdt6t+rZjQNTEChg+g9uoHfxb22CKo7nHV3VPpf7F8M
FTKjLWpiKfYLuxbNG+3G4OJ/d4234k6kK53ytyqenQNx8c3yBKzLwiC28B6wqTnR2tZnVWaObHrI
1VJgvIqvkw5RwA6EdFJGZLT2DAR78wiJYTDJLHhfL3YkrC/FYi3af8BJ5sW2xumeiXZgERNCsHU4
O/gFBtK+ql4N5HHXDXQTfjUQrnpv7P+NGERnSxcVvtab/+2mPK2tjK5w8QNI6Tr8+yC4RWJ604au
QJXgXJlDc7nqwpV/snriFx9e4xT402mkWKvL/e1gzrtnCP4pNvYWQz98BTPjxodvWLEI7fBQV2Hy
YK1M7SDZBkE2IHsHEM+bt5vhO9CwIfYWxaA+FxWhHs16XQPhVKuG6s3ImlJZxuf4b00Tf6iFXTIl
MM18qnlpx4+33GWkKz9Fd5LLaw/WuKjXBhgw/Y+Yg9UPHg3qIQUpiE6z5VqXfjUbKRLkC8DTwyvt
M8FGFpCfzabIEKs/EjivGpBNr9i5CQvRmmsjHsqb50GeDac0/z5c0nDVr8RZiCEUdHAgr/TpLMyf
WZUlbV5FmtyyfjwL/PKSK2Y3inr7ygw47Sl5s2KlzK7gS9T04HpZBmnbFK/ta6SPXmvqk+hkfO3Y
sJS24iVKsjrpyNPDRZGd89dz6tAou1dA2+3xGwhiFOl/BO4nn4R+IiVdtLWmO+XVJUACgTc19E7S
LRIH1qDLNqbv4AIjq+1LVwb+4RXwbh5yPCoIYR5DWBVlavpG1uv0bllxusV/XB7R/JUh4lvo4fqQ
eAu2FrAh3anyjfFjW75GammV4HfeA1f+62/47DED4BnP6HIX9zO9rgXzAJsC9N1DTqyYXUsc2aBy
/HBt1AdMCjwngQ/Z2tnyBcvyAxk2H2pPVw5QlksoB8Qi0h+B5+dZLaKH6f4zpqtzAoTipOMeR7Cf
nlXwHYaz/OVHR/pVBQfibU76DAgRre6ft4oUqXZXujEn51fRBScIFbLZUy+eNLhmG43RSA7Lr8T7
UOtIkZpuberatL4cMX10XkQqaVgIUfQohrYhUUy0NbRPxIxCWvKxdx+uetCAhIwz6F2ne+64bqaL
AJuZnPDH04EyjFDpHPex+qTxsVFQQmVJ5Fr+n/FAzwMrJDz/8xifyT4QEpfukoh66efjeKazMtMZ
Uylf3xoxsOd9NOVihoV3IePCqREwz+qsMJ6MyZlFLcluW3E0+Cpi0XcH6vgvp6WF9JwM5rJM6hcD
k2Cn+KFuYlz4TqB5qcYCrxprW0OK30+jYylLbjqiC3e6ZQ79QFz3zJYEUcDXu2ldU7u5Eump9EWM
UTF8+G67/aUyDPnOFThIiRDYYVv+mp7n2T/raZR+MRZPgw9LjWwwpkiwQL3Fp4jk+n+vaWOYPhqx
xgq/HCEL/+V6Ep6fRrCwatQtKPMiy2wF9bdNII2bBQrrH97/p+OK4982PhDf2Qas9I1HNItAQltL
zSQOInPNLQ42k8SzyNcMg+1GvqfwvMLOJrJrXyxD7TqI8YnCWkEuqyvwo61XO9HTGCjNdLs6bo6T
Yfg/VINeA8fsRHtVirBgCR3kXblYHfhNQqchTF5bl1tRKcptuXco4TxxRQSGfT4azL0U6qNs5jZj
RUd3oMqQnc2ETYpXRsSx8Da4UKiNPB47T+jXB9JeirFaWhhVr1K7ygrwpq1Jvr9PbZtEBgJSSOag
TvSTMNYhu5KInuulViTa9Wh2BASeQNm9gDeKDtQaED9/Jwh1M6QT28aDCSyg6d/z4nBV+ZsofN3G
iwvoCfp9cexByw1W5JO6zFy1aZlpeZxyd73nvCHGp+g1nYcZGxqcJCK0GBR1iXVz9AetjQ5whMl0
lA3Y5ymt7mSmT82gihHr5qBBa8+ss8xDKIEIncXg8lqrKBeMZC1COGTbhUipsY4DlYptxCGvgypt
FGMzXgZLboY5jgXnrOsBCha4SFApG5iWMbxMcrzMEszXUQ6DcK4zhcZdv6MdqebhDt8zSPeoQgPI
nFWG1rpbpi2FriuGJIs0y1c80506jwlqJ20py62hAb7kaBMNdSW9CGN2yBQjlGUdwfadB0rxQJ4J
1J2qWeH7lueuE4VXRXZqn1cglhZN0Eb3FXxbnYyfFTa4LumHHzJaZOVjkizwgLHHzPBbhChsChJU
/n2cnfCKQydnBDp7CYB/srwGbiWMEFqnzs0GvJ8g/XMSbvOWCC1JMlZdp8iLOOHsm9/SndeIlExU
l3pVdJevbRBSaAeZxN0jZXhY5vX/9jMl4c0cjXT8GbJwhd4mgWKI5PXxC9HMx+iefUbYMK1/JKgo
0By8BLOmXwes/L5l7bQ8KVI9kgYkHVDyeJzqt8+e/UHpuXt1IYzZpstMDGsG1n4S09cl9QPLmN13
VVfY8qtBaRslWP0OFzt2FReIncIAkjS82wP0hLCe12sHNQqPfJRKsJii2c9+fBVmEvaECDTnW6Gk
SmB8drnMv4zDe81fBY1FEhM7KsvTiKAQPVnW8igqbr3xhZwLexjW4MxPo/caw+BTTsiyQQJKog5A
M9gz2iAfqEOMuCl7gG3+bhSJ9fPfbZIqm0plVH+nI2OKprYDHhoCTyto534mjayvMuNe++H8hRfg
se5ZWJNyOHts4JCwceEn+Z6EkJNWs6octSInK7umDh3UgHMCTfgjtugdAy120VbfIFZv7Y+1nXWc
ew7E3ExjTZBZcfuhtDy0E7MkBnUvqY4bn5KXsFSSPkh99el7XPSc6R75SsI41k4FL+YszsrJT9Ss
QYLcAUC0v+B1TSDq9dkG8bEc9XynjYcDpY761w3pZP8nmyY2d3yhHeYa+CMZJv2TOUtl4Y5Wjsrr
xLY3a9EXylZ13vm4xQTLhq4ePiHXSD6ir1lZxOFzFXvwOwv8KR+/Uv6xZAc1bya/S5oD/c1W7NcE
1op/QZAwIJfPWi0My8jFjVu48Bf3T8s3wHbiUGg5hHetLJmo23eBIkwt7QZyxWOsFNKc+BAU4XHl
4E5e47Twfc1npMvatqoUnuHZFa1bRgC9K5dGvbAyGOZ7AGec8TjBQoBOBZ65TL/oENiKxmINKDOK
8wWnX08bal+0qTZkk3dKYWBrM3aEa3tXQoZK9ZC/PjAd62utuCVNmdnEnp1gg2fax12qvKOvjnB6
aY5wzWnnFdmzsl3a1X3sSgQliWa+CSsD18S9ejn90kFlVqCjSHeU5ZZlGnQebrN3AE/2hwm3Eu16
krO80ck1xN59MUol3RxblL/BjKtW9fvldZGIJx6l8tJs62lExbCDG9ynjRAQnzmq10Z486rGOqxL
CC3QuMsS60spmdgiOp9OM6fi4C4cXvC0k6maIefSnFkZelB1Bn9MGNAXO2891xqmVXCZH0B/aSxW
I3geGwJVc+Vl7uvrxytiBklZl/Q8IN90HG/NrEQZlatRaUwRO/3XpZIEDg1QXIQzMsi06iTG9F01
C6YVPKIZhkz4qWuDLp81b6huv8a9Lgv2LJqYw317pUnCK3uPAGMGRyVk5ggWPUNi/dynhU6EH55N
Y04sHnmXi9f1qgAlZ/ccdwtcEnnJbeJPr/UdZCr74egPzuZBXRUxvxXw8lya53jXK1XiUEK4cmKy
TLgqThT8TgRCl+KHUqZmcBMFv3IEsyQ338MGAjdvS8nQnDZeWEhTTkhWqP5q+TDkvbQ3KS/cNcIP
kRvVs64wIOhZx0d+VbhWtEnpwdokt4hMsWE1MSEy7WrsZCS/73w9DN9QL+KhbRt4fFDwf8g1FtFZ
kUQNlehwix2rZ53I30Pa+2TnPqtRugc7MpkuTp8OMnn2U5Pr1jXbfMIgJhamGeOW4zgJWuAl7nY5
6ShyXNURYY4cVRxSadHGVBzA/N9UsSLv9d4JgS/irsjlrP8ndegcvrjY0DarWEnKr/26N2cLWCZA
xTntGVdTAcrvBGqjp1G1hgD59LqGG33NcXrrFTjGKTaLZ+oVWsJb0/pJyl/3e4c+qNAvEh/49Jm7
u3HHZ5Any0vaz/5cTxVd47GGNbKTr7wS3wZLXjEyXL/Dv10G38kvuhu812cgywv9B9K9UiviMVz5
xxiBpayJ8gNk6QJAAzCiRnfwMCEFfAoFNWl9lajVaJUET/aTJVV6XiUw4uDBf9tWql5/oUn+S7/U
fe0DC6DaMdxjxyV7LfYRz2WTpBdfTyEp9ANLMSfZjnMp00dIEDZL3bYwr3Jyx3h/sMyjWlCYba3e
EiCjnF8CXzMCOLXQu1HWRw3NXpu0hBBQMo+5rJX6WrIQJj3GwwMQ4do4HALDY+7pZb/QJA34FMZq
LuhT7v6kyulNO77q+gLqKrqs2q14HNuY3Q58UVBBvlKtRqj2+BZ5T2TA0gsFwAAKQ4iyyVf2nPkE
6oQetSadpF3A+CGwPnIfPufQIbScTBsO85EHMPbzRNvAEc09qfehX1gz9yr+jTn+ONZ2FEThDKD6
RBEgaavz6r7Hd90yFy5z4MM5ec+I5rdJxUUxbpqVb6jveFwH3vOX6zRYB/x9XAoUmKK6nZq06GyL
8AjPxd4sxrfa7VhUH63IA5o8ozYQSLRTPSoCqKeCS6oAVzIgkq4DHMeIgRRSCjVfvJZaA8XMC17I
8RzbRS+AzMlQ3gmUVE6Akq4jZb453SeI6zhOchupF4Gu5FT1fOWbRxn/To9FbPm7TVf2ySs/IfC1
DY4VY2PeXvV3g1xqA7U1wrVu9mU7JHViUu+tJ9ZxsxX9N80AV4sMpbzX5VPasd1s4WkGEA9liJA3
xAa3SWVlKTpLcX8FM0ofIJ36XS7x2/Pjs9VJzEmd3yhzL3YAq94g3IevS3d6Ax6ou3eDCs0jDnHA
TOk2211F3nN4dOUaiDyKPYtO6dY1vCcsYnMmRlJYsSagIQMU0vgFXTAatkhttr1TLltPv4TfyJXw
JEPqXUaz+eGZAZAQy/njN+AgusDbhlEowTPTAsDd8vB7g15VSaef0wNPFigNWPygDwrorWZAyijQ
9TGCU++pJhVXqrP/TdYR/qWai2pItNs+k4AZ9ohWUwOT4QTFMpd0lTYIVCHbtvNbmLWMJdickBm2
DSS3J8mvJR3Nwb90B5pzrN0+MHneqv0Ty1FCFBTNhSNnXp3WgEOhF/0qy0TpJrUSO8Hp0ydXqtOA
Ky12nJUc+xQrAcgx6a1nSRH/OpILOn8PLPTgKgOKvNwv/qJTxP9xMxLPh3ENMIpYQUpKuQaX1dh7
f8t3IeWn3NV7YnIYTql9uYnPZ9ZDYywt62vhWUyZtM/OJRguzp1fhCg91LOu8QORpWEecd1OySlH
XsylyTTpnwYlW2yHIMxQmyfglOynwtG+MBghAGYaGXJ6noTeGdaMIiCyCq7mgcRPsrwzPcWa+T3h
vVW/WX+Ku1wUHBZNIDDdijTPMFIVmWhetclb0eIw5rCS++wsZ4rFnqfu3/lFXPR1/Gcvb81s/bLN
2OMqnf6Yth6k0MfP7UKA/m2+/lcpwjGWhSy5Ws6utlWzjNgEkRpmTMaKpLl7EjzBGVipnG1/DsZZ
l6eE2kkVtIjkNMNTPCG/YWRV9NWnlQ5r7TmedP+plAqf2Vxqz1EvXORpTqldN3dct4BNg7PEZdPd
g/64qyA4cGq192gQZIiNAUJWSOlfDpbcLJL6qm0EfavPZOLoFOz64AR/5jZB0m8MPp3Z01GKuOb6
Id43OVH227Nh9V2/IgaK9/3ZVl0NfbiFd8wqJUCOST9vJvKfN81DbQp+85qA34SQZmXzW6CvRJyE
5fs6myeIBVkhCZDiRBW19vwRCwrtwCDPy1B75U7hBoMnOyzB+DzwbTK2OAw8S3evD/FEiIZD9dGi
WInDaeEMjtPZn7O7MPxDvRUHTsl+0CBAGx2Zo4hYLbmTQXvB6zgUddWTJD6jgJLptvs6UlB7vxQP
JWT49Uoih4hceTeUqkkyL8OWAjIL2snjq8N9OZeqmtYRQaZevALZ+d7L6NKt6XC0Y2NfMH+jZX3o
sGsI/stHEz6KZgw1ZdrUdJ/p0HzidDSl+4XVipvObD8pZaDsDppTPXSe44/wgIVuLaIjJVY1yvpU
nuu+Y4RPxYifCVaAvyxEw7BNGmjDOpIb/7ONXMfHVl7RwztIK1MW5E7x2xRtjEeLBnBKKBsecywd
lHr495jZRl+wyK6DzwzTtMYzoOu291b276Wm6ZkEPaKh1UFsJA/giL2Mo1R6uluLkF9bJ9u74KVc
Ds3RN8WiRDLC4OjqvMHdJw2pNIAhr7/je6g2OgtO7WogxBU3x8qXOEmODnNA9kRj6UbENO+JO1WB
m/VTGtLBKGsRqJ4ZrnUtmEuTMPjD7/OGR08ZrBNIkA5rbSSacSD8WYG9yvpJqp9JsCYQuOSXVn1f
ec41IZlSQX4rjMrusoo2L0Ud/OmFHNWw3qtvXlRkoRP6uxW3+UZAF4EMn/TBsofiPFphglRLcIDW
AiGnYlWmNSg9lYBDxvzn0d4gCqdxyMaQH2FPFR660xU4gx626XMO2GQY0kGTGAEcMv95EoNkOYQp
G28s4SW6/xn0NVE+lqSqvAM+5gNiFEbJmvBrGUOmYNpWv00ujGpGiWCzVO1YV4y5vp3C98bZWiEB
vZ0SILZm+IxSvEyp7rABqgEeB4xLbOHDN3r24ZtJh5WnmuTtDVzMdpaWN7vU25XJAmUUwAD8MDyW
IndeZOjPai5XhoAlI+15+g950TIBFTkZnQuItLRl50jvGFOak4lJneISjVGdH0Pi/D/BWBkH2KYJ
SuDJesrFRgydylHWbwHxnbWcCfKxWwsMFdbM4OeWv3LCaieo0wYB/qDsF9EMO6GKiBWxJ+mvJtdx
vUpBhrS4WEsVv5LXclibznkA1ZkQvUGMwH1ROHJJa9SXMZ45q8OPaQcCCdSTk2LTA9INl9Xc+oe2
X5daMFPlCP+cP1lsLLK5jHrjL0ah6t6whLwPbUgoIPjqO6euFCqjHqx+H+eMGIXweGtTozp2B7l8
wPTKNgjIENh6KmeSfsC3sn1Pjp/9DdjO/Z9DttC6zQPfdC8a2ZD+/TM8FyWI5dxEsqGiRJA5fmfC
juFeQTxFcOUMrIkHkiI+ndvtF41pPygaVQ2CfjZIpnzEBgctxyDAl0yOMlCs2xBhA9iuYBdCpajL
vA3lPmMQ8w9pGfPx7fakfEOt4QTlDm+Q8TI2oQK3JaJGsVkFeS7D7/sChqMHoWqNisLHMxqY+6s3
HmfcUSVN/o8h+1Ua3bmnK1b4tPggqSSK4SNWSriL51Ut7eXbWFff8vEnW+N4vGx1wY52Rhfve62u
1tZkxdrcZ9wHpZEqMHXBYaQSaUaEEvtmulXmUaxbCEn0vNMtIq1tsdTGzpzxY8gQZOS/8tc+0WJN
dG0xPIUVZoKW1AoSoSLs4v8TRfAqlTQ78JN/Hpm/36T1TSKAGfCXl2Ff+ViPZMRxiuBlgyHGcZHR
wrpFnHqiC3mtxGg+RuFD6SJ/O06dLrF8IuiV4c7tO7Uj+PWT+HL0+j8K6MSG1+dzuIBThW018GDF
RWOgT1cxB66N7KQ94rzi9DH8IUiVKVXkoMgbBGTqRGnvCTRwy4T3z7B52RTZ3Uip0wCQBBdrgcDe
70sjzBopyZvpD0KObRMqCGmvlyTzPJAgCCJ8Bf5Cd+T2sTDC74H6SUkmflQHmKN5fVRled1zXp+a
QvnotT/1mw/vgRF3DoR+BBEq9QxDL6Q8Blmnzc135a9PVq3j9rce8gW5S575kOt+x8MniIDdSVFy
yJtEvEybDe2XUFa8pyg8FTISR85YnjO8eM4zo3i136t6T0sVNFgdt3O2yk1fsz9KhVsXKpCQzkLg
Xrhf7RS4jaHTBJyRmhSvWgFl49vJQN+EYLMzVdREqfOq+iRiqsD8k9Lbw/nFPpTtp+dSq33nIpCt
mGMohov31fh7+4/UrvYnS85ypBKELrsqLc/VRCBIrSDf3bIQETXkF3a+pvIixulPqxGfh0HcOPDA
W8257uiLdeypji6XBJLdFWD9O6Q9X2fK0faP7NfadlJ6z3lOalnP2NBBSrUB0FOB1083LdYYf1yy
nGPUUXtaDUP9qGATVYDjgnlf+zw/ksV96ReOHlfs/wInLopZRbHYerRuc4BkPJXqe1vZhBwcnPwh
UFwoGNLBhKVQtFrra8LAWRh0LDpkUID2Y6a4Tgam+JmRvh+0Lxn7z+s0prQfw98mR3NZA8hHaXrU
2zPgjI0/l4uGMSX+xmwGMG7zmWTQudk8ItOeqpOVcfKGVOM6dJCB36Z8g7WGc5nEwD5X6cgADz0j
9SaCAa9s7/wSlFaawCw7TsXs48xAo2WsB5JTswyMzvQaWy3OkOIvGm9cFIvAi0WzKRc6FPmgTSba
ICxrB1xnKWBMdmvLePGk4p4lwhwb0kZiEw+a4jq3C1wC1I/L9Wqrkv2wGlM7OtCaCSPiA/xAx2Xx
FMCxw48fE7PnyZdbzR9uKc/myfPXXGvqYY1epBdYIOV2AiwyZw/1KzUTzNBaMXIxuVgYq3UsIxhT
c6ba41LoBlp69pJaZn6smJUCxLavaD8TBak5ZBqtJo5lkr54ZMe36R5y7SXDxeckOzhVWL/Bbusv
GufAfnTVqplmnVgu2/ZiBg0PpHeON4Q75HjkUgTPDaFH44P+0dPodaLwfUAKipX7CiZTk++GnYOK
SZnIiIAgdJTN0E1rSmbxbdUlGEaX9bSvK0DiFWK+66K+7r13qqtQ6Ul5CL1hG2EHhUX2FlNMq5rw
ftJi0BHhu/A33fNZ7fhrLqdGj7e/SB2ABEZ393kbchcd5FUH1bZmzxOkmLegdqUTEVGgRlTXx7rS
NCS4gB/KcIag33I13uoEN9K7Og/Bxjtu2yajmXUuKKbL+G/dJ9JU/tvVdTQgVBfQ4RbSYPJWmrGz
LGRfOULqDulNUPukeJ4VKYgIBmU9LG8x1W2Sr+NHLKqjq9/i646wn+ERddtPmXGXMTk10RZV2ydz
sB8cb3qxBw9/7TNiHKyZ0MuMD2YvHjd9MeK/flEM9FXmYJLCL2HWj7UdCi0tqR/Dj9Jskvs2+N0e
/Zx+CsuaXVAkLdMnWWwUH9ehMkazjNEHLvbNXdR1PKWdWxFdDAXyj8duHVjQtAya4E6BmDomwYLL
BkKbVnkver7Z4K1YcJiaTdCskQsg8SvqIoze0Dtdgsp+5SocOb4CFeDRXFEvqmI/G+GOqbmhWWYT
I9ECXjXaJ03XtAHxlqGSlcKEB1ZAnOj641K30xpBa5OHTYDASY0mgtB8XZn74E08NThSCkqqGS+E
HLCKtCWeXAf3/Bw3qauSvLiA3m2ZJVkHsthQWEUcNJ/W/l9/WOXo5wV6cGYY6aThWGaV0daWRNT0
hJDddu0l+wGsItpcJ15VJK6Yu2juO1XGYBZfKCdVQoRsdhyYRjZezilqj5rLPfi1XEMeDdd71dlT
vX1c/7w85zaG13UdjY8svlj26EXbq1cpSH8cgvYAPW+K4/1QGct9CfKR5MKGBCZVdIe8X8o0EczS
CHjJrnxs+cPGizCiCHHwtsxi2nSbOIJw4YOBM/TUd7Vw9UBBZHVYG+st664zWrONB6y0mNas8uy0
pRzqNfXerqC6ys5FJcDlgqx6NWPL0YXrsFaqDPPqtpJzWv1z9fsroL/Q8CySrr37LtQCO88WuTfW
IAfMsxqCoSaBERTegwjyUmXuXbfW0ool0R/64nlPj21rEzeNuG0P1Aei/MHtt5DsV16BHVOQrBcQ
zToK0Loh7hj7pPBv3CWs4xRQqOIkdqV3/0CeD4v+jQIRnmQwQ3uiFQy4FoCWcq3v68Qft8d9UvUu
lAI5sx1+t9dUfsNyamT6bTupvUlzxrC4JKHwHZcQpkLIWGirFzeyQtsbqVoWxLfDD/gpQi7lcsqs
2BkkEQu08ulZpQx+7I3uYdSXwiiIV6mDZydEhlPFs2/Q3yH4lNOdOyIOXIMIe79JpGlt0Q0Vnnum
qe+HMhDyUNAtuM1EuehkdqWV9KGVioFgv2XXl1shV9xbhZeDlRa69+bdYssTOQiUa5ruvapN16VL
hCkkpvRBy0yEMBTi2+4Lxv78W85lpaC3pbDJeRIFRktEU1GQYlcaVuqgg0NmlDzvvsfwwYe9sD2b
fvwToIlzZ26s76dF3m1vzmzqFdpfynbiBpUdfz5R/9xKyiMMuH86jwOeNKpcF3j7MpqHGIk1u8CP
Lrv/Uu7fWXcFfT3ycDFwLz6APYx5LNjjwtL7zLA6liBHoOKLzrlwa9gPEjNZ5Osk3geQtN2Yzqpm
F8p2LuEl7TifGYtPdDKenuoyJQNkw7pqZhQKpV9pioo6myXXMerOnRpa5QkGhyyFV4OWKua6iphL
3bbrn9JdWWOmVezdJ3H7ZuZjkGuqw5I19GntorIngl3qGaZuiE7bxcaOu2nO+CWQ1p4mawGIfrpU
Wm0HvMYW9CFYujQMh/eg4MP4d3+rhtztGFTAJAF4lWVLfh87D1o8L9+Bf/AdIz4PgQrmypEcCkvr
tKrXKWINZl5GzWfy+09GUU1deQVP3jAGbmNTXSXoM8hVZ7F9VV7IJvsQx9yduWZKIXo5Go4WldMH
7yXGJ2ueXkSKh/7u40b20ZlbDeHJgztiodT08GsRe0VV3+MM2diz4MhPqQudvu9EdRU9UizPHTsE
q/Ugj6Cxxu/4jHFAKqz4pO9BF9zAubO0W6jJRMnr5tJAOa/LAVOCoT1ZWEXfABGxfrt1kHkxsbJl
sVm0MqIr4jocFnpY4x/eY/EIHzyAxml9iCTj6ss2FiagIdeTuq7kWOd5M+w/tgT/ftBIYmkeYKqL
WfACVnvt3HBmmJ5JE4CO4po8D1qTrWm1g7xrIaUYX+Edu51OQtejQH5uJe5LL8qf+dYL3DxTnFcY
18YnmZMQwpAyCUjdosKsXmPM3tgaD1PHuWSrphDyksuDlqXzrb3Vk+1qkqCV1GIwTDbfegbdNoAp
dXdNvo7QsubPwO1CyqEG1YDQd1G7BExtpL1/4oVGlq3jGaEmOxk9atc08C9gx950hgbV6GJAvpRW
XAk7e3Cwh2+QL7K72ENZzDUhb0KsB6BrF0quUFrZ9GBiB92ZQuFB3+gYgvSM9Ewz0ftmHrp7pI1v
oSGHeG0zzT+w/5OEHGM2+W+wSduEBm8kjxf0oANY1CQriiawTUFtFEv6xwGEWuYQ/WaP/cuIPJgI
v1iEQ579E5iXAxNLQx1MlvDCM3ywE3XxK9hGBr2Un8shbfzGAn+O5jTg2su5wyJ0ycsS5oej5AGY
cO4uxW23h+FJkRmC0gXgo3fyU+Z25j5DGVoXfR5x4/G/PvJuQBrGxOiqt4ZmNookKnc9fruE1H/p
8WESXF5PNwbazq4JjbNcVOfJbwQZ1CfZcvoqZus6VCio8b0Is4tpAJG83Nyr25u+siJB39NGJcL6
p0hvUSGIej52WetM49gAMjSsh+SQM7AoyLVbkyWcM+9eGc4tZdOE23loAZAeElGHjzDuMpP32fLp
/YeI6Xb8Jof2Yik0Sz9GZ4H3FH1HurcB0qi2GAzYPMMYWw0IvmEzsXv32Q8aX//iKp1fkKOTb+/E
UYJQA5piwcaaIf8pdY6EMGe6Qk5DvuAHQAsBiK49iVVkNal4jEol0cn9UeA5GbkOaeboXCehlrBC
Cokr+tyLZVQYUj9+mjxxG7jkyYu5rGIbJbxXU4rlOzN7EOV1xf4V/ZA2wwmadMvm5spf3JIAb1eA
B30+Cq9wLZfDhCyC9gPjS3WJKGd62V3YTvc32QaYgXcMU9FIHeQ6SnkS+23Klo/lZHCHp1BRwVuQ
ouvx9C2kZ8QvJO6dITm/N+y95fUm2DNggzy6c4qN+qk5MLu+tnWXEoKZUxk1AcwHlJW/hJmn9ibR
h25uTPfzbDwrZdxZh2nCOcNbNupucLUkbovqe5fiG6mZewgPkYeWehxfmRvkSIHjQ76RJJMYaEPO
k93yrPiCBbypw+AOapXLrYyzQf+uU34KvV9EIF8uUvJm5Vg/dFcC5ZI3qOgyhUqZyQ43u/e4GZ/k
3ifwviYqcIxkuQdfGY0kQU/MlN8GIAb4I3SIyFIuTHwCvqbGmAPuPf7Mnn3rpsPFm7yTRtLhBo2e
zKHZuGdpuEZSHgD32zxpc5IlsMZaI4TzFl5nSLAcQPsN0Hlqm2txqaudag07PqaYo2fCz8Kkipek
tAeTd7X4R/YKm5lve8VLVZXXj5XglWnIaEt5i/CU7sQsmWEcOYZKRicMY4vpMYNghiykGmOC5sCA
E8TRNyash1PXp9Gykn/ZrJq0rGx1Ds9IPfwyMaSkyrHUJFnsymsdtO9mTGkHqUbnjBwkmTrLliPQ
UgiX/LBwDkzpiXAAOLQjsqBvSwHIAAId4PHc5oPNISh2T4iDfp8KGsCPNrRVdnDC6MXeeJqjACaP
0bb2e3zcYR6pGmUtFKegu5SF6EqKLbMtPfq7VOpr+I4p8py1rXUQE0dy6FDJgSflR4Teyx7Nuzzr
VKfZjWFWnJhbSPRP4hqgm0aAeht9dvkYNhxLJCK2gDe2dFENgrt9/mKTgeGruIuev9wbdCbtnSPn
PXfA1qfgotpsoHngBX42EpYBY2UMx8V1FDRzob+Uokimf3HPrQZFJtUF7LiVcQ8YOQXYz5KPKazO
+Ht16MoTSfXpW6otfLsAk1JAkPb0Nmq72i3ZAhPXSLeUr+ujnm9AJZrMKmVvHvbcEZd0INRE/auK
uLMLUeLAWFga2VwAlUPRWQWTvjlMBle/RB+35V7OjrpdQxQD2H7w17IsQPOl+to2yRAdOTUC732N
vI3ys2tl7a/ur0fb2LKEe65y5yoDAgRUb7tYz664wCsIPZiIKhmWGGq/ftMhlPJN0Xnf86gwXMMy
xxIzfuHVmh+viqDDX/Ovwv+DO89Cqhy6VySJpOCnnCt8GjMGwmZQ3dk9Gs/bcpbcH4dyS7h3hYP9
erRxR5vw4RzYf0M4KwTMlCWdbgPMaKq0J83VTl1pfT+AuT6Pm9PDMJDk4yI4c0ynHe3RuG9CnwNo
szjOQjneuLFqXRKWU4jDK2cg8hfJD7Rrv/RjvSZJlmvUPOSAVtIRtm/90VuM07Av07bWxvMvRzaq
vHmxPpJM6pyJjzpFc4oxvj1rWhTo6QmWVBGC43dyiYKtP8EzvYvoDRX1Y7diuAwIU2o5ohMeizH7
ucOOKCII7MrZrSh4N9kztNzVFoaAioYNnbLWXoMYX3fmA06hZYF/LQR6d7x/btjKDIJNo427LCqh
zQdpa973JITan9qWlXqwPuy6h/EY/dv7KbOkJFEQXLTxZnNsw8ZyDPRFq5AeYXqNenU7VDw5YBrm
DZAgkVzD/rK+AJSk703l3wHIZete/Y/1mdvMb4y50RH4FCsXY5tq34S2qf5wq8CC8h393Lql6pYI
ZOamsWt5Kq4s/nRUPwUq7JXSa3A2wBVtDoQLjpFJ6u+0MubJVOsvNp7IWuv37kKewrJx7bKUie72
IgzjzQlvNcpM8YueltCSpF6BuuT62V79ufds/UDKXgS6GvsFRzPWuoC4pD2SFHFcOP1XMZecbnrU
f1uXr/5NZS9TvVEtFrRvgb2DNSeYd9AF8NZHVX4jPx4yBCLDCjmZk+5T+3PqC3hRYdrH7xXRrqmI
tVR0zTgOmYLCJKqi1zNaugBMqoJDmKWSeq5QeldAM7ImRcO1pHvivH3LsjkA/iVWPYpNEQNdDIEV
Mq+2NJO3TyU1GZs+bFOaxDFSoBO7bP8qQV59ujhgLQ3qQsuWEcNdmhPKtS+/ONMSUef1CnENx4h9
IMB5JPVhD7wyk0vupxYLzftDCGg5Ba+DUifQCXQH9ESd9W+uJNgHqhQx0Orrdhi6u/OFvUzlVbl+
FB08GuJ41U91r0TshALcIMBDMuIWezib2swFwwFJK9GYrRrI0RMWZz5JZGSHzHKlpItqUFEpTr0C
5rproQfNNfOTyQ3U5qqbqMI4mZXiKMMtBTBVhShnee6UBNSoib7fPdRgik0CtNDAC8yowzKCvu3l
rhOanQY7FjTWz55wTgbUyBGs6Mg0xvltyRoqoQJLD+utC0f8BhbNYhkkKyV6/aKFEQBFvMUUcJG1
af4sc2T3r/m7dQhbvOg9jtiQBHJy5SYlzrJaZ4/37coLqVFWcTCXNOHIoBNxMWrL+aDOi60lywQn
ZSfgWuTq6UZfOdJvTQREKhGTIxXPTQ8CZdPenYaYhgpVNsAILYXg3gNeFopNzvHO/JUBv1BABwUr
ch0A6m5V/WO2WpLl/l9e6PXaj4DlgrxsCZFylnK12n81bk8d9zv0yJUCSVmJ+sKGnjdZGDjkv/UK
voEhxhcEcjQnlckGDmovVmcmSuPsKbkIej9tzids8KdTdQGy+wTUrEgEf9dJ3E9RaeU1JzGlUnS4
f7mcFvovHrMj54/Ci9kBk6AiDSvEQKUHHEef6aPqYBF4q5stLZWuPZYJ8AA78NnDpu5PJh62n8pK
7H20fEEZAr2GdpqAyoI2bHFQaEZ8ETWbItDuFE6M7YgOl6kPhQ/MnaKObeCGi6ChrlgzUizi6Os8
N/KFXKZ26lX6pi9mkZVib5KpuScIQJ2GDHU1sGWpdV1Eq8xCK+Xs2YohGUyhh12LMiy4bdgVrAvs
BSK+shDv2/NBYnIIfu6feP9dfe0ZnKarlFCB4/iX612lfTRu/mppx4S25ND/0X+5Ysh+tNlfH8pJ
UfxKp1IgTpYpIzfa2H7qIRizMLq4SsHELhdbUDvBdYKiya39y7s1SVAJMXP08fuLh2dYtpVtF2Fx
9c11qTxBDpw8qtBjqBKH3Gr++W4mTIenU41xd6v7rZGjBgwYUg60ULPqTUT9DU5QxkpLNakej1l4
08vglDv5AdUwwG6DzooUTOG2DeNxhjXCAdHgpMKu4Cn5ikQuuboXgeSQQlOTQ/bh5Q7xMvPkOsX/
cPRn5XzN7ak3yTl/kuuK06urqYKtisDn7H5JEv7rkToRsH3quXnOdyx/XQ0SWv8wMEyKHURqf4ym
O5d0SdD5BTlKFAGhLUbp/sB/9uTWaQZPddex9UkUZJhQuxHBnTvh9/MMjLdLLipg80ktSsgDNqvi
CterzD6PZKUFWIGM9H4oO9sXXNfLt5VD/B+APz/nUO4hJeBkqAkZq2TcQgPURzCVv7UddE1yni+H
aGc7ZjfXZiw6seMxr/gzYPdbOA1xwJbHglpO1Q1oHzN3GWGcubmGeKWXvJL6Sa0qgCq8RGr/XrpB
k5hrSj0e4Wcbxz7s0XOy6YGciCIgtb3dr5ZfAq17qU7AWCBr/XFHPqL6AQtllacvAxoGOa+kzbiV
X4zmbQefIuZhu1ObKgZ7xVRfx+zQPD76mMEaoId7PR+UCi04gEq4H+1PK8dN+mSPuxdN5md2Jqv0
IUybmnK+bB0WBXkUclvvuKQUFk29Fl+Esf+IDQ0vWQE7Ku23+XPvzePAalEXayVtNTl5tCklveq4
rdbHjFnmnNCJREF/nBQkgPuSSFchS0SU/d9zw2gFBROd5qDit6nzRHYzSbjg0iUoWQDz+jQCoe72
AKThOEVQy+JLN5/3/iSQnH6QzMG2cXgSkO5/M/MQptjwUnQeqfyK70vsTe+Z/hwuzCHDC+PhbOF4
4geJ4zo5FbGTJNbPXgQOBKJjgXbEzFrQb6ktNj0AUFNrF9bk7ZeIs14AcM2u9TmAc/MgC8bcPmLb
GfZa0CpKXVEFAj/ezw/7wWBl6fPeBNBygTBiNeLs5C6WvSDHouEuZ0OENTBWNgWSwe/D6mTJdJ6q
vM11cG08QT8li4k2o2N/fuYGWGQiFv5tRC5/+88C9lunfN7hSi24qjECoW/FjQXMzQP0H2GPVnt2
5UAmjyKDcGd+7/2skvsVwMfryrST8VMgztGHSH8OyklKtlk5ro347uDUSENnZQPhPizDScx/D2mU
naQcdOXVyOU+Go32Q9bhzY3T34ZFFdqxvMsrDN8iQ6jRAa0KYEpCHuu49ypWAGMvNKlbgf1YZr8x
jDAbRCw4EoCO33uMZP8srSQEiv6K05w2EBVu7hRcXnraqYImRBEaKXHwf9mWTyufFFmf7GM/EPua
uk+Tf56B5kweozusZrZvqYt4ByElALwALdiPEvihkiCzlmsuMrUFRxS/vXX9ixKagdg8vujCdHNM
hocc1yiKgxK4RiE+oWEPZdQhvSQPKY6zWTQpy0l3YQPvoxL0V+GCoZ3cZHT4jb1/Xx4CV30FNxP6
ZejeaMLbe8Q04fs0WN4JWh0kHk9OxPA28nsYNJKrlMqBtpSwOKU7xl2ZYkoLKRNAghQry/6zDZb8
rblIQ7J/SVLbe5ZZC4pum8jHvSBKeb0iN7tR1W1vwdfWRNE0z+frKAzDHutjM8bFb1Vs2zoGHj+S
I85saoWrwZ+v7mYcWjJPPZM7PPRocgr6gfbN57pmejFGxvbJ82+wiXcD6OFkhv4VLgrYPIZR60/0
Im4wvwkFNCiX6hTt3RfbWMdoxPXpJmmlfLC3IglrCt8fej/tbOr+9j5bvb+0lEEBfuldAviX/4DN
ETrKkybo0f54vJp4bjeh8mweM4yDmw6PhPCCnd5jAyNw6riatzoXQT1LOmubeQ0NLSk3bvfNkBdL
7G32qdCsakyXxFsPJr88zFDfURgURS7x4RGD9A6oYpbSFbxGazCFz2A3ZzHR/83SeW7BncAiUUHa
nNEPSezSOxW+moTLd+UyNaoNR67jhuZ7G95cciLnwwDONCakCC/vdhzslaVNC8C9bT+dqgXdo5LM
wrssn/PZitzC4s3oNs2OBhPfqQdIC2uCVFNJq6PTByIZZM1CES2liSIabxJWRn+56OESsbBSkAEM
vgAlzZesRZcSyaEIDGLtl9+y4bDxSKjg6aSgPHzaGaaMGWsujCFaXGTP2OUZKYbqvxyds3NTLQvr
l1SXa5ZP+N/912djV9xjIRxOst9yb4VtOx5eUBqJ6D6bOFXobLXub1M6uL5fZklc1Ug/sF2uzTkz
H9J8oMEl2sjC1VBteTRb/yf0tUMssAGwKFmmwNfO1wdVW6qHwNrgLaM7xwK2DN8wW//cJTOQTFWc
n9DxlYE4gVsyc/FiRW0VDvwhBgzbDRozMjE1E66gVfC2EM9QY92HWQThIV7AFOcjXDiHDlsL+ifS
shZtCS61GOwsl6AXz63kQN2wJ1BJt3LIDHx83FUyrPG9/aBLwySd49xvXCsKssMUJ+Ae7TI5K2zM
kMRPd1E6HbMJ1mVOeVUJaRpEXUD5MtPp54D4Jtb94891pX3XyxoziX9s+cNRGf8kb0if5uqZNwZP
OCUCbiyjDnTvKbeupgkOYhh4mmmRbo5JcDlHNeN5Pjz7s+VqYFPh+p3m2FbSx0CLgv3kHESH/qU8
JVe5EvTKaFCFITjUcQAI024ryEb9HUs21Dd+pLFJhBiBuxlGRUFFLyrUILJj33VbhhXu3OKXxPNS
D8BmRTH8GJKtu55OVNOt0VZ3MhrCrUCXHURQj7F7eB5XAllqZ4H38T7kY5LuibItve9OhrsPEZjz
XDd5wEOmWWGuIirhjXdpNUs2jP9ZDbEDE+cm20us09exCgLolw8/JKKIwFP5Ctmi/9TVrwCUx1EH
rI1sWEIgRekOsvMkL8rjmjFCM5+85uoAutjeEvbPsQ9wWdgk56H0DxXiPcY+QYVnNCtSf+L8N2Ub
YsMNmLR/gx1isnH4T35jox2kUtrdI39H4irY8VFei14qZDiakSZtZOl1afDXgRIMBqOr2ppUeXsl
xA35gBsMRSfpbR94AeHOggk5a/bkezMZ85Sgj9JBZb6zcv08dXrxAA2CSQbqljmvqxHHnA+lLKcL
SN6xhVeAPu5Q7VqFcvf4J2W07ulmqksHqCURcs5E+2yZeSmJpsymqIRJOmpm9+Oz+w6EOOV81LQo
048uBgp8a/4Zom44adG/vHtAmvKu+TRBeduHiSyYzheRQWJTA419NgCaGVr1FJzlkxXVGHCS3SWa
QhTDl+1sRWAnowghZWvPiSzAklR/SdQT8NJJtJe/6SrJkgPTorNgq2Bm9jqhqnxu/4ZeMfJVMlOw
3Hq0gwWNr4+TCxTVMNCYy+fIeSt+GjF2W4AMafEHDkGbqtSPsV5h5jHEdX7aey5NFcU8skkax/KL
xUKJ4VEjUrSLD0twWTZ6eEImEVpa61ebP3xryYqPMQK8uyVM1o6pKGtfC8GvtuVe0BCQXNKAGITY
vDBbz3FzucDvbPiljxcPZzsbDXTXQ3HQF54KXeBK8BoCTnyWjvMLMdFDoyYT/xYLNIlGncYQSW2E
9frv75SsxiZB6E9MdixCoTOUCDCYc752dPD29bHLtO2WXPqrplJ5trQ2Y5skBko0qeVjo2xd/a2r
YbFz8Z9JBehgvDCnQH9OPYu18WoVhihTNAI65bD0CAhvoVXPl70ufm22973HLWEv/vnrJV91qq+y
F2GlwYt5cs6o2xU4zFs1fH7xMilguIaBCVh5HgkOrPslMx++hz4IL5Nfa5NTT1ZQVYoJDyud/Piu
DeTVAZL4fN9FbNfo7pLr2jqLCxtGy9VKcoBdHeK+oz8OAYDV2omyoQYtPtkFFC7wyIWfD0dhWJKW
2Gh28po5JnIoZf3XXZPGD5eXeG69KtPbY4qqh4iD72uSVj38aL+HpY3fXm7ntWl74lEKPgKwLGYH
0B4QQGhmE8gUZItM6Va9W+4l9RTFi1HcbB2EdBHioDYvH/EoZcOTeDy3mk6JDnjY+3OtdoB5BjWl
oxLc3IOa2NT/f2PpAbBBqgMAS2aDne+ScuWC7BmIwoMxL0t/L2KSNTv1rdhHDGzRGzP0nD/0/Zfj
qdCP+Zzr9RiQtDsP2XcMQUPrZ0WaiD8ubg1Q87JvD1zkhgxELau5eK9qfoDzQIP+0J29aRwrisDn
3COzN4s+/u3o9x5CmtdoIHrtnmeMf71Zhwa7RkmYw7uZv9WMZugbpz0y8JE6LszSoSreXldTEeGJ
V6btB62X6pXzYLcBDwBGK89SfivUrtpPofLkgzPF0M8gxOZb611ZNwhNxmp1/AZCyRKkDJYFUaiQ
TnZWbM+irguRDv82w/JswXYXRzybGoQNdGQawLK34zyDddvLIKrUupFjn6RjbA9TlP2zRh4vgDvV
CxmfXMH9CxfTRcGqCi+Yy+pnbChyMSAPXz+PvteZgW0kC0VoGGX68PtwqF1N38/5NbIq19xNW5zG
v8VVdd0V8Fc70nuCz9r05WZNkg1wBsW1vPNTX/xLGt+BtJcPGuCLMCLXa1jBid/2RODNoBLA2Z1F
Ih7t8euiaFfP8ha3r9QPPkhkj8P9Vosrt0k5iEK7jy/Hvr8paumJQgmqO3W9rfQOukpx1XgbntVX
q9YcZqabCKMSqS2Ae8x4+j3bgNDihY8kT22m9MkB8x6lMltqWMOOVD1CZl3ZvsnGiJcLAJnMrGrV
NruFdf2B0I7U0VxXAbaDnGCm2XOQ/MbgRF6rk4OxrEaUzqmH01Ers15CsBae33XvuHeK36DGxZ3G
8Vvs4r5uN0VdGZJlyrqHjOOaUj9DMqEbSD0MhOrjO08tEoSIqqcYFuMLeLdGWsEgwvvDvSEbDWgS
2lxzH7GTIGyYnkpi9G0pfdiCBgGVssBVGzdHNDFoSJKfTyIXZidfH9RY1xoHoNK5fLNXRoc/GwaH
uKyJWn18gg3S0KJhksd0oUj+Thk3zehWQQC235yQXnWIe1KqzYKDv+I/P+1gf25ZJIWGnHnyR0nQ
irolzQd2QoxYlIfToRO+MPFWtqZzrbkCR0EuVW9zhkTFxUzKJ5W2ZfeO3EU3y7aaFH+fKeuRmJ1K
2F7GFtzCdoB4I7SWPIKAxtk3bpD8CpJMuT4x925pr3oKSYjcn/rAihk4YJll86AtMP/3l1Mh4/4m
KJmUDZZkrC6KtLRJjWGfaeQJ8cskP6ZYjj3uNr5LbEDKvtNXlJd3ArulufvRSmi4X0JYMI9eLL3J
pW6YCzpCc7S8k15uGdIHLynAvO/V/hEPOO3LsFqyxOOLNyQ9VJGEtD72RxWrnL5K4nSGOxzelHtt
GmKirWkg2d9vju67EhaemYN1BhOuXjJPbJ6bPBCeyI+04zeKg8cP7yhb2FJXCMduWpQxz7BlVY9+
IE6OzJPf78TB+dcdSqfBwgrfgNXkf1ZNJQlmCfzocg1wk5ExAuPcGCEaUIF5jHyWB9ye6toYyxpy
a0eJ3KEh8r3znsdFfMhgbeKT5nHTzQ3TWAscQayv6QbjNOeoKXdphhadZ2hNmbgEHEwytRdUchxS
DJugHC5Y873OyccLuAnkfGZyLB3EdfLQ6hCHl82yRujsfHfameBZ9HZccazaOHbbHNNFWWc4ts4V
qwpJ+zmi+PMxRfBcgumfwV8441d4eRYbpt4mWoywOTC34BwzTrj2k1waUflrcFJ1ksLTN+NK1usM
Cv/e5G04FQginQNl0XcDq9fnoDbdag097+w8XF9fRNE/7b0qpJRoKK3RVZ06Yoq7OdAe/ztfUPIn
yZduYCq49UR0yoafTUJz+gO8lFjf0HJp1VGen0TotkLOQ3yN5NmpdeLHsHKYmZaoe3kV7XVkxANP
4tYsSE34zJmVSIUvgp2RZ8UQdncgPl0y1BeLSukoqpxDcQ9taxhyAZCcWEor8W42uXfP1KVnVmrm
LMsiiXpwbPOkzXKPj3iAVyL1srBVc2X2viYi0rWDgjEulHNmHLSbnHpcqtFI1YRw2nihp4eDLRCu
5kTISDsKicCQYDj39AOXZg517JSgjyhXxKLZPPeqd7s+I5gzs9/eUmb4Cup58IEsrVstGF08j8Zn
reesDCgP3Sn8x+UULW6Wg7dCbR9SjcRqJ9t0HvKv0pJoGizE+p97wMrFU2z3Pt9WQoaMc/3VJYfT
ymDIr/1SJWBWJs0UFgsoSGN1KDC0wmXtkr/LxjoFJWZpo5qUlsICh+fI8T7EeTqmebrHTheG/6Uc
tYIwXuav0/+C2Lc5h/kSB4AkeCQefgtuXwDTymulBF1MZTUFVIop+8AoosPda96hIbAX7hidBU9w
/r1kw+tyLp1d29LD2ryb1fGlcu9SxBYB/arN+uzpnnvBmTHY/TzzEY+kwxj+9+4GzElVE35ePTiS
DixM3YhY1/f0WFmk7HF3Xp+TkTg2U6Fa7kWZ6PlsTACRHfRE3R6+c5aCirw0wEPImFRD/Zld4b8w
Vs2N+QfHUboc5EEdufEDaRc2mIiHgJtdbLwYgxptBeQsN3m20H2sFDkiNii1lHrTOIXIJn3uG8QU
6FAB9uU/tUo0n+oHQZUhOpCQ6pgXB+PNQk2ZqmJhAGkM9wfOKqlRyD2OKyvw/PIb4rZgGcBr2VPH
y5cMv3gmC0TaKKjWN8iGEipROFwxNKYE85qEmTEQmU9Tt17yD7FpkIr793K4k3THB9aT6lwn2C1+
KwCSozFakUqxJagL9V7FoV2Siwhmz8gtFXoPrNr+BDMzKooB9JpA5TkohSFhdxYvJDZlqeDGPjKc
3ESqjW5LytzzjaV1nMsqHD/OzJJHGgJjbMHRG1c26I+rmbArPQNFKTXrAlDuukoqeVwrJS9pmK/a
uMKnmImeH72nWlF8ue7VaW+WIHiCu44lgVBJOonuMLsSeEPvyIH4bpoPLYarVLKUixzO/jDy6m1A
g5DbYtXMjwGg3247aGXO6TgL4x4n9MbI++KgeRdn0x5xmAbxk3OqvrN+W3T0nJvIasYtOXh0hb9I
y4uBwvSAVvb8Fwqa4RYh/sa656iQmI8caIAEbPrxDjQT555kWb68I1v4GM/SLvlhiYs9FV0ud6Og
nR+YNdoKI1mJ/GuH3RbAlHNJlsVaUTUytLO0ku++5a/dfb6StlOCXO/BUKhs0M/HlagHE7IwqGfG
2nOoGtKy7OCbnO6Bmc+VPbITM0ubc82WB817rcSEiBe/qNrdjt1gOPouA5Xo5uHPbIwbtaohkERg
NNlQsxd4AevsWC1ATS/aQmBEGVJ9Dq7VfgMqt9+3adCT3RGKIGBYQNww//53mtdhEc6nU78nXeEi
L8Kgw9+9jraScoZMWFfLysHJtePbY+784a6hB9JQuaPpDPW3V+4/RgPPIKKC21A0ZSSn9MvBo+8N
elHiaOgMDV3K5qayjzbqFI8N2JZWp1p0BDyh4eVBZE08vDkbotaL7EgPQA+0Fs5WSvN0H3rK5t8h
nNSFcAHKfcWLbUFtJjsBlN9llPio1WAGVI7Oeu4+DLeJ6Ks1PHitjlkJnd1s6pAjg3iIvuDluPXZ
G5YP+v9cKHPapQQn3In49bAgWhvXzbFXAzUggipWWkyavXcViR1kd4CWpJIzaQpzFNwqHlVkfEte
OzdO1TLp0+O8cc1pyXB6w/dYlBrflecnqxtyQgmw1bwbM8mLV9hhRru5Z9dwxHV+hF/WSwLZjb2q
QUxqaUSAaSLzkwCVKmYJUj+IzRjPWKCptIUOOLLZC5Er4I5hU8pt8vjDy84oAvRar7eGicoCA7Vr
1mUeib3CkJ5RWIZMBOoSCWNLNGUjmErRiDvd/neE/IwHwM03Odi+yjd6lNKH0bIsfEzUMlvc805I
bjdYT9p2qZF02KYZCiT3VaZvW1VhfT1Jj56zP2DLgpfMRhlrRwVAODdKQf2VIoBK0iDsSFGQP5R5
5y0VXXtqKgcuDH29IX/LARZRXy1gK+oYK5+ueurWSVaNCPKPNHuyXMYd+FcSLo9FpFjgYvg1HqR9
4M/Xo38jDinC8FhJ4o+L+NOIrY97U9llhq0KUBPX0k+FVQnK+U1AvYxNeC5LAon8wbAVkR3s1sJJ
mxhwL5B77zHYLD9dXVA1SE/pcaX85slALEJhDRKGVRPMqMy2BiRGNcND5MhHRsAQsoqrEx8FfEb0
kBElrr+K2zvumFJ0vZp4KNpEBlOMhVq4/XQxtbngEbxU/DRXJGKcILoeBVOk/ibRwcBQRrMR9RzF
HZaw6ArBLzBTq/Aq8iweYCtqrgyG7Fc5ShsLzXLU6rQXEp891XpASusWbrJg2T4FYuCrbrN5z2pu
V+6HRLOQLYJweesAOZkO6avWbO0pkicem7gN4P44kc5k/sPhOyVUNvbkTK7YUWpm+WTzMfl++Ghh
kV39d0tfSDj3eXvKnICeedPDxVldgFwdvpKlyf6MGoXeQYsTjVSVDITJtHuGknOHFFzUg9Oe1zjk
TEt8E/InYk/Z5ZDW6to6V1A962KTJfhyrHrMdJ4i76K9PVPa4cfEw5ZbyOQKSv7tUbfeAUoC3bo0
VOPESvuMUf+hsGOh/53Vn/OSLJI75lStWHGbqmVWtpgKzaowwXteFSuVGrUAAoJlBNfG9tI4KH6x
F8VUxybBcYobZUSpwZkdQI6L0on2NEfc5/8w/KLK8+fNs5o4psbcmtdcl6sFiCr0/wa39FEdXgep
BvS5sqHIF+tnAmQ5qVgGPO04KDk+WR5rXFQe7t7NoGu7klYhwuvNg10Vl1wFZKl/D1P4SgdRiEsA
Ky3bQZUN13N1P/Bl8xqTROurVXlg9CObnJMkUwjbbuE/6puuNNyPidoJAUqmQFk5CUpcBfbhkrup
IjFcHws6QFF7fE11YF8ijlz16+mSb4AgBCSPsvg/rB8qIqi0X4XuVYxoan6z+uIzQGf+mGzOR8lf
qWss8rIYlma6mVg9tVR4eDgaviUE0Omw9i/UI9lRRFT7uwcDiInYJqmSgvhQgQksMVEuC4PEXYUM
v1Dd1vCvxpL5V0l6Bi05r9AhPcixV9/rn8Tr4ewTKg5ggRFNNjvPTUlGd1aByLdnzxvjkPCMqGu9
HwjWp7JjjbJlLAgpyFg+hQH2Yl0m6D2Wu8cEGsp8v4uYywX1WwZPOgbbgOMo3k4+A6dOJgVeJvr3
qtrdaK5XUG1+15BGnuxnGcc/V5Rp5yuFcn5IwS7fqcxxAu0cCg2eB+7qZ8ewkklML6aZdbNwEKjj
PM5yy11K0sAVN1HymbbD987FipbDvvSasmqmCBwKq3sO6Px76xd788nw8DKKGhw6hV2TzCIGVGwF
DqOYWl28banMVL750rhsZkhkh0CnzVURNmmKyyuEa7LbWZ5NBlizQBD3nRsyTD/xaewhZp7Ex355
a9osYU46GqAmhwukh80CjltP71LlA6x6cPVJZ2PLQiz2XcZFhLOJ/FORuhVsb7kbtMfiXTkWwRZJ
Xv9uE+tX1K3bbeWXvB7TA3ljp6rpMZPLowbPB4saqeHBACc6k6VRAi6l1pPpENGwKHvHWVlx9HKe
i9ai1QR3xJB2xLx3hy5UkMw9Y2/yKPiTR/moY3Ym6xb6i7ii00fzSbOe2/SAgacAIUo+4HHa4v5g
lK9S8SIOCPPe/O8WVEYejLipqU1oKiNNkFt+p7KyFbOVpOCL3YWVDQ1d/zrtu9XXd8HYb6CwrBKL
2a+kXfx29hKCQrDYtvw9RhFL8X8KuAUWfa+6yjyo7iQhyO1bgkbRjBkx7Vx41UIkZfLoNvAr2xzP
ZgarfkYXyh+rQHOQdvZGPYBTUiQH7HVgAHl69+pt/WD/9hG5KJ5eBo37fFrHkkrTJ9ro5aJFnFMW
kB6BnXkER96J5a3Z/v3+wXZQ+yGYNUwCgldYk/GaTyEeJ/ggE1rJfS37vPSvMe5ITqyDTfrgB1DP
zC+9VCubSjmn1P3jCmtikcJ+XfVHL0lJpODW9MOR0EzYfvvDOREGoZiK7P9vsaCLEI7YflYg8HQy
HXqF4J/MhanxO2d+Ux8GWz5s8q4AzsSa4txNW6NiZI7l79Li3MEka0Rk27QNYHAS3kGgu7w4nVKj
4GoxZYmKfCr5X2D1ke+HcVdlfSZ8YECoV9cmX/SZAeKtvYa7GSSLa8dk74+YeFSAJvC0cQh5jidi
UyqrJF54KF98emqf2Wfj1U9sZJzjZoMLJg6lCuHdZeHIyF1k8t/wwY/K4axUexNbsoZDyFQxFjUO
D6gSTjEs28MjyNQyHXz/mxsvHzpN8l2O+KaDv3g7N9yK9YXjEmyVZTxTdTGHm99zgIMV8M/TbYrP
REMcDZT+vrangXDRxH6vA21ZDFpWmLwtRb8OPbqfrmBSFXY85IGRtGhgTCaa+/0Aq8XfvsmK20dz
QzTqdRpb6vDgeGOxpWLwG34eL+O2UEqFsd9cm5RF9ClGuhArvJIUgsxCZBKaay6MN99W1nVtz6Oj
+M3wU26izgDaw7okGWbBswC868KJWmqTNzT73uOW47Md3CInCO5vGGsn2wgfsLbSUtNgB8qJXF8r
SB1lwjjxOePzPnOQ3sxk+AJ/k+bwqTPNsa/3ihf+KnR2EPDQm9IMkvzMymyGYYR855a1Qz2Q8GlZ
QKx6c6JF8E8C30sPc9dzvN5fNqs/efqssoI8hgvwFnCL3R766t4z0x8/qePs6vQr2C5HvqDgz4i4
pTGzuMGYClp71tVjlUUgX6ZEUGMMXQ2ND4iXvYg0sswk/e/UUYA9RSsKMf0g9wu8K8CvS33e+X2Z
aC/gDrJCM0MT63bU8+gtzf6ydSgs6/Qs7O8QZmwlfUDNxxDaliCNSQ43++7cTpk9jUXDrf2UUK+M
YasWimyQq6o+VEq/7kNTRiEK33aKQV0VYrXXnaryGObOCHBP0kaAXM8O/cJCZm6EsiKmG34YvB/U
fmoVrW/5zwv7IJhTyqRyVzEtZSH6hIMxhR3LwtaB2wZtnKywrBWPS2JW2/QN50WgmmV/BONas51S
9nTyYuv42d0y8ABGuGFMo6jCDXx8Rm4GApeo3x6hIYe0YKHVk9U1PZmUP9Fufc+CUJ8F8rBYIWyW
xY7zfw+KueLszUVrR0SX7imfXiNhaj1GFlGlBtMxju5bpujfiwMNUp0EF/xeLSEdqqIApUy6+8TX
ofTiKMNZ9CjE9r4EwS7qMIY4CUMh43YDV9SnaQ2vPXNd4Qc3VGMmtqEd4bToKaH89T9N0qkdJLUO
e3U8ZMGAUG9juwDVdTHXqOKYFGV+JU+dcg6NkV7AvyIWdni0621wjYfN9qcGg6RKFxp1Uz60RZFO
2qwQO6AuaUvMcMLELuO/rVu5uqi6YWDWepsjS4U/fgvgnDxSYbnXtlZQQGvU0vix9uPMSk+mecV7
jq54RZPW0jER8M7LEFQKC33sFWduizZszMyKixLfF1aSReM5Uwn6n90jp00ITQBIppzoorvOOnV+
poeJ2o1uDCy771LsR2RRmClYADffKa4Wd9nQPm5GfNn29mJJs9up/vuAdIy/3nopChbaDzv0wN+L
ce29Nh8DanR/rE4ORRgYVHk5jTCHLRBdDeA8i97oIX+NWmedn5GsvW2PiTZOmNsaege1jpOtYsMm
uUonPiU2+BsTDAVbn0Uuuxuj8wf+AgHisSzPlA+kgSU869K7HC2BCqjt9wc/Go/xbOluaMgyqXze
5wbyHOKkQdADWwyHKP0a9bl7CM+wP3q04IQgXAAIFUA9SCQa/KzzadqibovB3ebfE/CFbR2dVewE
PTQCT+TSykoHhac4lhRuJCH39ZXka9xl2CxXLbGhOZT83C6qGgMsaIW1eHV2mY0XwAlc6bAvNuiI
/1ITcJCf5CObVEwyjO6IEpG+TogrZcayrdhwjqJqZ3e3shXyqy8hsOh4Cyp/86LAKvKjgFS+oJjN
r7ilusoEhDars1xc423tmYYrXJM8UC2g0CRrOxYUUyIBQb1l8tqnYetBZWq9FViH3vFy0sINX7u2
HLuS13qNEo4DCs8qbtfy5/xFOykB51Wu2XH1Kw7pdRKzynAnjZ8aRJspj25k1Ks7CwBriR00imot
uvorOWJ+8LPrRAPJg02K8/DWZ2+WR6TFJvbtad+jyhm5qwwuHEQtb8rMdGjwav9VqrSniDANkrbb
jWOHCT01+Kr17I9QmXShVUaJpnMqZJ8nwEaTv6ewkN5NaqeLcLC9/GYkR8D86V/QoJq4z1TN9AHG
+6/LYIn6goGh4bhs7TjjNhmoSsoMDN3e062kwYWqnJd5n+EDmNHU3RMsvLzP3P0tPEI7S8sgDIp9
IcGB1vfv96+d+DbESbdUf9+jWzmz2CebmYDVFgpN+39xVRSYPbvVn3FoxMPm3NSf/htaEW8LGscL
dI6Xb0dumonkRryRvqZzA9zLTAzd+KHYMcpfw1oWJsgfC8ru8zKAHcaY5nBrgza5eF/8O9/g911o
l3YbHxK8ZjCmM3vzbaK1bnoQBD4vKnBYSuz0DCtbNhnnNFvTttJBhENHuvdkavOi4ujjL63778/B
P/GXdwwyfst4dZeSxaThytAU7QhTozzth54XYZSHIjZMTD+1r2RjlSp9VJeV55eupYkTVKAUazSM
zhrJk6jjISJSh8Nsn/sC6tVs5cYgH7teCAuiE1uZp9dCK3gZEsk136jAbth+9GUnzJNR+sUjj3fX
Q90n7uTn/LQ/jgrhkEQhq4w0jVqXH6wi2uwvtpHQFCBXUtxCrqsZbkcAxCgszRsX+GtQIV5ZV5st
FXH4et9FfC6BZY2Bi2ElDVrzXJ5IHvPSHbNCAVqwGcnMlTNw49TXGonOdA7GTIZxWNRT3iwh7b3i
zAFUVhNbao6nq5NPKnsPx9iN/9e5Hq3cvtAIoB0mDiOZ1hM2L+0eVfqc57ycrFB41j3ruaQNVpkA
/Wwp28RVkt/vF2KfSpvOlIT0YcSWjv4WvDOiqo/vWl9pWN1GHoo1P9AveIG6jxFWCKepwCQyTdaW
W31JMIwnQPbPTMxHIc1lyfaYgLwFekZEq70W4qJ4v/txw5ZQ/4fJ+iE6zDlnG6nIYI1xAGbAHqNA
LIyFIn4nK3/JE4XL7ksk3Yg/OPThImAT7UlJ/9pOg2zGPIoNsdZNiL37FV3qrTnUkz+WAYjTMURa
3V0zfoZZWGiEA3bpuBw2Bhc8A2n1Cq8mRKINGyvIT6IUPriIckrXDlzTYbAfaoXIUrbDhhZUlen9
OFNbwyUE+JujJBw/34a/GHP49ZO1e8L9u9qdygAyBiUOZU7z1nRbVShlY1mu80WD7/29Upm6czrv
0xgQyQ8Vr2nuJSyM64PxPC3Inpv1bsBtx+woCS0DHymDbtAgDEHaD2/x4VjrVpCyzRFdU0iwCrNf
8YQuG0IP3buCV4sxmkqdBcbmps0MPq6zZdp1E9rrwSbnF/aoTaSVkVe3hXK5qbDVDr/88pSFwh3B
noITCaROLymZNwYjlnAssipitNZXcwxW++tVqsUaRHQbFQsjhG+JuytZshG/GmQCAMd6mWuS/0GQ
XMNTGmzWhqVMnnQCzA7NFTtcnV3vD5UV1EyDSoLv2tz7y/DeWm9ZhfHbggODAwKX7wsHBbtGbzdh
ZgedbP0eYDCQB5yZNdCiRdoemWDpWRnKWDZ+CHTXgpem4pp8V/U0QbKO03VfiXI0/wyC8+/nslPC
iRTb/5PqablWo2N5mhMR04tL9qtoM2hhfReRDSUZzVW6HpXjAtSVm5LnPyyXJk7gJHj/ur5I/P8V
CMDGuGB3ALmHRkGW9FZ9HRT8ttMla82GjZMihfsFzImJ+zFftr+UiYfcOxxkxqVhP7oQ/hkm/YHp
lGKQXtCvBqnL4uaaoiTOujq2HdYgNj0zu0SFJvKfxdNJX494B0aST/e7aMnn0zLqf9laSfBZ5h81
WuGt74BMaiY+5P4myPbMQtQ+ZyAPmD91+0vb2JMtkRuieDgcirD7DiJC2KZtcvqrjYfS2PREf3VR
53rChi/vPXyrYLrUQYWEeXwZecMi9nMe3Ub+bhdNEjrpIB7FfKXKAG4hucoF6YndqccePBkUrb1S
N6r6JgAjyW9C+iCtbh0IwOeuFPOjGo7GaGlyqGFeyk/I6Qok8npSj0b3eiWj85I1TWrYYtHXSiw8
gTnB28PN7B9VXljtGK0y26c1cok9QWmPYDIYQhbIJyoIZ9+Vq79n04jyPUz1Gl/QICx4VC6Ap9Ef
RCjKLpg1J34JS5mNuNnMt+EQYQVK+GCtvNTP9EV0yy1a5+gLCuLp27ZPaTqxOmQrhEh+J3Tpge5I
BGrZ2JHDTBr5naiGacmXf/+7exIQxrwZ9Noy036eQFUgKBKDqOBDeZ82H00rjXvW4TbO9QAU9YJ5
yWu+bw+wfjVLyMyRcsQ9k9qtCH6OISVJIZiAKqs7t+D4DhykcIm2jVBycg5TTdVhx2EdsZC0SESA
N1jgCfUM7rHVtaoN8Epl5cRZRUNK2Bq624aJuOcexz7NlgmTH9bOR+Ko/fkZfJJg54bYA7YGrKGE
whtQf8qH/j4soTZJ5h6rjYEbvFRRW0UM7sjg3BmE6nXIOkXkkotpFSpNhBio/2A10fJiUbFcx59N
5sQBvn6/5YkH4g0Sdow1EdXGNHBlsv8XtqHYy9BXhlOXuwhcxKvrT/rZpfrd0xcC7lutZEOvXjWv
ZDhe4Bigt4szZQMdz147vW6MnvoG3a8j1VswCAsIafvvAHyb97uETj3/L2A65Hk5WFuNisX19Qgl
i20bRmtfLpouXRp53yEZsaRB9fwaGRItKnXdOHCBUip/V9rJMouT8qo6wS6hbhK2Bkr36XWls5op
7/1VmNJ8pnxln7Jnb2UGKNPNpvun/dX5ikwygO8aSyOd7MApIGZAdg4zIyVOGNOhQn3M1+TtrSHW
De0ptKGdR7sa4VDZfTdaqL2Y8VB3ddorxENqzHNPudgSIjzINbI5P/rGyhcTnn8K0x5bJJiI/V81
qGaDh1lO2j2U+YDQjM+fs+WJTO5aj1BgE1ZBYNrTzMrBCm8dsCkrnWe9X6t3606pJiJ3KwFVt6R4
4wmjeAsKAGFgfPsofjHZFgfqunW3MC+vfdYgBi+hmoh7ecdEYPFcczkEYQy1JZLDQGHBOALZSZDN
ne/qHbnjS3j96+eEdhGOHlEFRXX9d/kSFW8BkndCfqWMmqoH7wdM3iMKTZcXqF2YRPTRmpzK6A5M
7FuS6yFnT0LI7Cp9s7f6trtUKrIcm0/F02Zl3653qClgFxqp6P37b3fyCuPV6zSnggiFkB+rYgt7
Q4hm9x9f3gt8mouCniKYa8+gt0ab48HhHWM4wXPqAegYzquVpUmqN3xQzqMs721sBId7zFwjgBVX
l9ZbB6cqs2kg3deidOH6dEfFJOqLgWPq7ICmwnkGyqsPehwBHJaIxdnRI4EoXYmOSn7SuU3hTICC
IoLOEKtUlNXj3BiiXnL+fXK75FMazSiz7Yc4xUkUM298uAcfK0Kn74wSYtFMnmAFlD2SxHBjL1/H
XxqNnR3DCd41rbm5ysBvQuapdgP80ILlZAsxWrFGssWuWY1GgCHM5CBygOXXr9+IdtFFb/tbF/cC
nHuV2pnX+OtQLLsDmKzcGLtDY/QNwiX1Uw2cThb5g80+Clp8uqNi6cTrYKbu9J40HZdrLsA6FoZn
FL5ykNfrOl4HAHAv4LWmuBiL7x2KGbYIFyCtnSNaYMlRji6JtKpeofMGoJxqIfvz05aqaOr6DQDh
oD/tPANUS94fdi15IgWP2ncE2QgE0Rq9iIYYRSmKTLCxIItbUWKLLbSsqT1gVVlExNr3HeR3GIPM
hT+J0K9Z1JRAykKjy2VF88zjpC5YoNL0CwNJVYWSQ0Ljpb62UAoGeBlcyZ/3asDDaovTB+JbY4XN
VBMCEYeoYrFhFRNazZqMCFEOM6ZyMMLvQxXGElPIFbJbzD3CtIyljr/TEUzPQw9iyoxf1vVcpm6z
HSSOVwghY08ZdgRN1R+JjwEHpnN0WUcnCNdcw2aZbsY25p08KPBOCqvjAfHwblEV0MbMuFbBkNiM
5VgBaK1HBukBVfC99b1WYW7iMORORFYPWGAYvWMACon7XCU/Me6GYkN+xkCGWnqm4gwZXpwmBo56
UeKDu7p1ETcpMXQVdUebSkDSEjvSG1SvBpSQotnc6ggNKAaoqepzRgRdQgQj4+xSLEofjLVbVM5P
f96GFkHgLzvlfGeTnBxJl8cpaR/8ouBpGwywY/jghgK8+HPb/SzohQyzOc9rH75UI1frpre4Rfnx
//D3hRF18rDTNiG3u0Vebvhvw6Vy1ThpRMqcTYeyBuQ1r/IpZJZxn7g35j1PPo3Xr/P/2yJeRFTT
/wo7EcQ4OSywwD11YhB5HjogpLVZwKFvf/1Q3rDcru8oIuUEGxS3T283SUxTCSJmHy5Wt6Sbb24V
/prcXdPyieDmwqbphvI0VWI4ueF4/0zASvPJ0aR1enAocByOlyWZJu/brUOIqUKpUwCGKT2S7+EO
bqH631sxqpIczEv1OCjqnqPAya5E1wkM8jPefIf1lhBykqrtSSOtsphfBFTnuLPrUO6z+X+8/L0X
wZOeStnCCyymsbvVvNgIwcYOM2bUfjbo7b0jZlPPgosCN2Xz+ME26WU274qntcLF+SWCEpAJUW66
l4OPQ2X5V8RTj2+L+UkXYnBBArLwur6AkggX75ml/oaNeULovyPwHL+oolFDEma4jRSu3y0Ba4yF
lLWDVi5IYQdy8s8kvAew4+ak75pEvWBntNfeW9lQvR17JXptJuM+2oiRp8PZjvLS8ta2dF2hkUK8
8pDb3UddIE2YAcc0lIq0ZLE3DBamSvr1Kj2hc0R9+pk0uuxKYtn60HMzQHhaicojfux2DgIY2Sjt
wtIStV0wZaLgkUjlwKJNBhOG4dhA3XgHxRDDLo6lvZn58lWYcZg+el5W10CENMjSLEQNojcTXP1F
w8jzO2Qp2/UzVhSxSq4++D0flNTYQcZu8/r7o6IOOG7jKmYdhFJejfMSKo8f3FNBdAA7+qVVLOSo
IFi48GTms89mRSc1XouGtEU8Q9NKMod2vBIoZ62qF1vDzL+Z8cv+lNpDzermonAloylIxftc5jpg
Lwl0NUaTK0+0AHZfnfJ29e9e4+GC6UdtACBqtm3yJg/nhqi+CHr40XwHpaYt1jiLv/5E8sqdcGGR
AlCNbD/BXVRxSvWHn3I1zaT/4ttayX49khbTeHlxTNR0+SvDqADraZ3xSIWaO3tCFa8oGdgfGWZ8
QhryzBsgN+tdestO2vGpoEndPgys6hufpZjoYTtJychfp2XcGhNRUVOfqi+uZaOot1F6mQ6humf7
C6H8LVrKYWiYM6ThKdEwvP+wxwqjWal2aA16pbcjazYL6HPH2UmuJtM5kg+TGrLP4RtgrM8NHDUE
wFG26zzhPhj7CB+qRL/6A+So8v+gMK0Asnb4QeFIunrMhIWH/30+0KyptkzKpXWRopvw4LXM6aPs
cTfibrez9ksBShtELhwiwudswm+4eF7L3GZ32geF+40EfD8XiISFRXsDT4HQGTu/1/T9fbl4A/dh
z4Bgl1LIGlov2fis1BVShG52XtTnIpJH0/eVCCAY6Oe1U9QC0Xxsa0gmIZIMC2Sq8pAkjQTbxdfZ
wLancjtbByEYgQvx0ZC/1a277IPg3negzLy7Iz3hdfoFZNiBg3jYcoBMc0XIsA+gt1o3eb1aqGdF
3rXWXXlyWYxD7MGlKI1Nx0lSdRpnPWqB6SZlgxBbVvTkRkim/+4kvbIV2AfofKafZ8nXlLlvcROZ
gI0CRih+0I9TCSHN15D9IWf3gPyDRWPM2T0pRGjyOxO7wNNMoFVj9E+m3w34++pCX3/T4n5coVnk
vlvtilKCjKY0YFpgBP3i9ja6MAgUfnmz9IbmkjURjwN/NYgVwmqpCz7WXntQyw3lBNJTH8Dm7pmf
yvi8dThlGhkVutDnSA/6NORGn0yPfeFJ68qckt+yjcG568NA3T7x4JPNyBh28CvX0wQTjZveCNPt
JRLKansXBmny7DE5mGSnp/Uv9qNCW6y6SG7LKUj0A3SBHV24dGyloiXHmhAco4oNM+CpizgiMSFs
xN9o02NXwsHQEllfzPHOFSRjw0pFqWK/j5XQjjx1lBB/mskbu60q0wF79ZeutdZ30Hsp0ySeFiJp
UjoBd++LtqQL+ohbS3v06NqVDgHy1VT3UyQKF4P157TzfhO6OCuk9KTTOdw16W8XJe1ZHuX0c2WY
uRhtouH+JV53LDONz2IvcYX4NA6rtodqHVE1LzfuBMypndZ88raIq/UvtZZKXYF72CQuaGuBbN97
IwPhvvsQ6SeEp9zM6zQXA7c9j659IUKiinTWizfZH6wwLYdmUYRmkuCRd9GzCpUw8zO1QuUeDR5n
+qt6gI3YG5qJG6TEmbC1UWBf2FyyzVOokNe80jKMFrTkFdCPMpWEWUvl7NH4J3Z1pRMZD3zpeK6m
tQQo3t1c5PK8mYJYGHenkF4gjd4CxTYgNeAlqCNcn2kN7vD7Pwb++JuER8fdVp82bp+twF7xRZbR
VnnFblCPaVHvb8ijoG/2yFfRclyP4RwE/rLV9AKRY59U6RDryCU7MoV4jvAJkcGebLvnfIbLAtVT
fh6BNW83Jlgfv+oL1s3QTg720bGywZRb9S0MclcvHxLlHxWNYSqpqMFXA32Yw/5Zz8AVvzUmFlSi
hPg7BrsNOhiCSfZX605tokhNwir8DDecWZEBTA7MzAXJ890fUOmd3urTFsEcJpbZRp7uUlABvlxE
TUO0huEBh02SmLZOo3NcXi1mrof5oYdojMJPvYiCnTVcQ5QmCqG2Na32gxdxoj23rEU5dpjWB8ND
ktALfBAyRNl9Qkb51gnIfO/vaAjKP5knIY0ZRfk2pWsoqcY/VmE6ScC+87kvco8RvWzzMwTuPUTF
t+JfvWR8f6R8IopsDSPvnYJHoPRMVWs2+cApvGPoTbTqLQ7DJ0AOdwjGYX+z/4oZs9a74K1wYv+r
l3LkfalzSdW7mkS1AlG3L6tP6Bzg1cIZs3oLZ5jgtxeZ5PItagdPi9YvR/PWOerA4iM2SmOd6Qv3
2mt0Hb6XRonen0z5nPcxG1k1+KMmFQEp/FV/SacyJ3wzy+Z0Al23FrP7YT2N7qoztVxp/9mF5CqF
uVTiu8AfGFP52v2rlil9VrCixcth3NujKEI8xEBjpp9dvOLKo2hDYjV8xWYXDGDaMJU0Iw9rBUzZ
BzM1+k9lWH90riUqmcj62eeBuqUDegtzKLmRk3u51w+3rZXfswVZi5HaVk4HeuJGccMUYnlJ56js
1NljhhwGLVDQCZoKB9mppcByz8AZoU+DhkFrEJkOPSmlkIM03S2i13d0R3Cq5wPyRh0OyO7KPcvj
2aNpRf76zbNgNQ0goC/RlRQ/0mWsWrKKbMIse+Vi7MVRCacCpfR21rew2nICTGzC/WXhWGt51F7s
v1DBphmnUlTOkxxIILlBkbauH3v6rtI0O2KAb5z3xfgNmqSBmZ6CKz3pxaMr8cWCrCh9HUBtnqSF
DWBE7T6iLXZfSSOM5GIe6xPqRWxEG5ES2TrZImK5y10IUepE5TtztWnWo21LE6vy/E4lrnKac9c7
/+2wq2ivZkO2XCFgIdzVo4bdnW6dXmpvBBiZsWUdP5fJiaA0EL3kj6yY9HZNyg7j6K+Qj9D3EkSO
36X7o0iggFS0OhjY4JvfNhtKG0bCygRDR0WL+WVcz6fAkSRYBlU/RbLqR/kIfB7nNStkhv+CknBk
H5umKuvDa07TUtLOiUeZ/xX+aN/kCz/ZHfVRdg4miQmgTsdoEsae7RjPUwvDpuxvs6w4QERVne1A
wR53XOUc7j+WQldKK9xu3HhUDAqOkG1d5gIx82Hsz7vAU09ZOIzOQAoCHApIfYHavH22Y8fRbpTV
Fa5/GJKGfUdXWAiUTSbfJlkLRX064SMqDdaYsFCYEZuIlmOpgRC3tkIELVW4lmnKrmDRlQswBR7f
V/gUwdIvloy/YuTSuFMJoPhaRLuVCAxU9sSwkVjeBkdHAFGTsjBR7ZVrdyojWaqaKtjSR0al9ALG
17Ikxmhpn6itKfs6KAID1XcN4+jyexuPk/R7px2rc6e0mV4LlEDgQMv922FqtnJbnHicxkCxNWb2
LXgZbXpnbrcKdMOX3tbJ0kqmZRg60urpMUUgDp0Y86eOGR3UB/FtUuaFh2lr0UfsW07FV35TsjJT
VX96/6uO7QV0RbruVpwpy5C48afOI/v9Yb/8Bjk/vao5mbSJ9W2ERN0b7rbDMoRAZ/RUCCc5LXE0
S4R24n5AcsOxqvwmphLmCtspqbLidGx6e1bl9bkKvEuANOMQTMAF6ZXxEjO+aeE4rlYz+awx2zPA
jCQnaXdRpPzMQ7NsFSNp44G7pdfJxboxTqZHHHgRy16vZ4+dxO4XPHtdPT5GIe0YdkTdy3k5WR9V
Yr14I3PMwA8p723Stp0Jxp7bIeNQHnTPu22suKwx56wbOJ10cTltxc3vuK3wn7BNTci6BbsS3H+M
4XUOVPXQiK2LuKezjFvoY7CTAyTpYJxLmWZo0OVhJCzRJHAeSSvAnJqGmrywZ1hgg6bh0K7ELLSx
vh1nHSAohu3FhtX4N6VKDQUVA9AHxsJI1k4jbyjbWWYXjq/dL9155LFrzv/t05V4lDUXPqib5IpD
0KKa6GoyLbwC9RJirZ6p4y9xGdQtU1sXjM1dP9aHNhKQxPSYM88bXdvBn8VI9jzpkCyoiwvjvFvW
Yg2S41qCLQ0L4NT/7uvs7sNaSg43AZrmnKWB5Ocr5jZBkep7pVjZVixSrFnENLWuGdOPnnmLn4ze
JBSg73oNXPKU5Z09/R7h6BBv7zGhPb3UfEYx0W25/foKwuxaebuYabMwyBoapi60Qi8Zh+xFXAjX
oxQC6rRtL0KUQqH3VfeddtoRJvNDPzJ9Nh8ueT88ekO6AEuicH4hojh8KrDwxtJek2tDWt3CvvWE
VZoSGS9XXfNvmTMTKGJMBS6QIkiPIx4YRDC+HokHWCtdCxDb3to07dRJLAuX+Yh905SPCKfvmB1X
iR7AB3ETAcwcOXFXp6AQySKwS/P5H1K+P3m2imZZ3ZxsepdOhbwh2gexrLbdHJjAj+Q7WwK7npgq
PwdnHxRBlv9irDXPXCen8jeJGzqm4zKW7jozqdhoVTY8GP9qEML0/eDTTI63jsyP+7KKNVKHBSxN
r+shqkuvoi8JS8ZSo0NRLEQ6GQK25TCR64HchqLfBE9VJSkrFze5jlKXcu8PpHy5W/ITSCzCcHdk
OGlBju2lcQDBkb3SVrgMr1HPNbas6U1VEhoqMsMcaaAPmCPN9xxRylrxxZTVcUKz1hUhthbYCqXG
aKS9FXHrwdiSs9SDjgKmt/wfLIJHpC9W2ebj3/tN7sAe3tTLOy0cKxTjagzZlba3WFEWbtmzL0VF
k5T2559NWlG8BRtSS5Ahax5djZWBGOy+lMo92XBfUurNdRVxs2716UxpmdFHciqetQ5rF/mjKcRM
YevZT96n3BeANS3d2UWUdQfOuVFEaoDzPwd+PPHgRtWLJnI+8t2IoThuFDWRSvrDkPe+z4HxE0br
hkATz70wu/n8t9rz/UKjiUYiesf4Rqv8OYnv61tkguzZO11bPgjDPycafW+IIP+WwKEWbm+/gJcr
sTrV32CpvELZobHQGhMjjvc9QHwY4es60EmTgueY62LHz2XXiIeKqgOmXwoDQipeVQPO2Ztb0dXk
Ess7sagctfQV7xNYe4khZ3OR3ZmEKtU7BHjqVXDqvZCx8ZShuNSgRTUTSlViz/uMSEV8OWluNd5a
NqjlBZsgzOsbRNPqIaJapnwZGfPBAlU3NUiHix+pgJqPJUZHvoInpbKzSQ+IXLLU8u3gVSK6yAum
+neIZWnwUCWBQz+wG3OAbPeKHyDroheTtTejMHApPIYZ/G9htDHpAxPd6eElsVJIjMz7TOU0Nz7h
wqcM4t9zs4RLdpi6iVkS3iWpgX/aWINjETW4xHlVbpfKKCf7lvK1nQZN0uvEtfUeL8uh0xsu20Yj
5df5fw2INclxOjk0Ejgd5yDnWd9GD8TbyDJVvc9ludza6WUdvmsLRbEaDfXD/GLxbtpp6B3rcLfa
8/2fN/9HY+ajCZW5nVSpLKJv9HJoz5K5OetMcz+imdyrRc+HLPvfOI861scr9PDmYzqvrfcxuEJg
NAjkgWny8YZO2hxJQ/H9w5higD6WqceLYm6EpCqBShLMFWCzpu5dcPN07+4hkJYuLK5gh9wiU4Yi
D7Enyjvyc83KX45cJVLso+1Q4YyOBphhYRDIuy3MZIgm5JIcith7Fb1iDRGmjHqq/oBg7HUAcvEL
g0Uyvzj/UFiM6i1U4xZlmtCwfECbruSKi3slXPhdYd0DeOiyWfX+0AxutBmScY27cTa6S13MEp2x
7bNLA19MEasB7G6Yeori9kS3CR86iWbKRu5gldsucX1SzBr4JyrcUNPNvMiZtryozvVnXySaksRn
ngaPt4dyRPlPfEkMKEpaK3oZq3/2KiObLh+Pfl8cI5HqurXLKODrYH/bYJx1VMfmQK1nc7PWk2mq
hGp350Z6EcPWp2tZ8m4YWxEMTCjiFy6rrxTdAU0srHFVl6a/t8xwHOW/Ts2Rbnd1BLMNrY0eEqH0
QfOg8SxlOWMx7vG3LxMDc+8goeFk5N+7NVLI3NDnukIKVWPSwUoHuLrENGheIQ8Iu6WEAtoDHZW/
P9pF458t2knj07sLudvUnPnlDdtvF9RChDVVHn0f9NowS+ACmyu+CG9Sw6YFa9xQN2D1+VzMhO3k
Wr0JU4fkyVXBSakUPu0nCvZo6WhB668g7A+or+y27F/A4P7yjGORgp7XCBZxugTzS8wq6pPyMLUv
2TrPTynkiKZvq5imTjCEJ1u+RLR/N+aJWV8qGJTqHdvjSG/xdXOeQYa5ppUfX89CAp4oKU1+2idf
bpW0t4C8zFyeKhbg54PTi+1BbnnyAjswgK9egYH1LhR8ytIBeN9KyLQRpqF1vNCI213Imu7zV5CA
md5wvXE8h1nzeZswX/F4rsV6B0U7/Q7XFySFLgtv697H0opstJlVdfmXsOh0dXncAvjixbr9fdh9
WVDDzLzqKWUVrlxmtbgIppOVgw36y/Q2EP1+qBWh2JLnzjzPa1zfNNPrXPAFtRojc0d5GPKv+G7g
lMepYt+SFzTiZV0WsJdqWeLtMby6p/gxX0GentrPPCIqmgD+jrBWZh0u8TRY2SftdRZb00KnA3U9
xtVB52bmmjj8IYVlRdYm9y7fWSKtucijT8FD0lNBF0VCR5mP53KMvm8QYYRWF4EL1Zd53GmfNd5h
TckjfUxNY2zvy307BGYLJU+oEEUK6masDkyXHopoga1QhmuBNV5pSPjDE6/yBOQ9klpq0mqKEWyh
5KnMIQDd5NU8LnXhrJo4+D9WLJEU7IXHFcUbdXaX+xMayBCYDFBFBc9RHgynC1eGX3GSTpPGcRtU
5DKGjlCJ+ioK1PTVAjtlFMtqAbJzHehK7RpKdleG8y3zaJa3AuOtKfJFuGtBDyKwKPLvtw4zIVMG
lbhiRLCoKrr55bQ+3bKDCuZ+QxvvSkpD/njWlQ55gSUGMY/XIv1mVgOxZH07IQzR/sD44BGdIUa7
e8Qv0/nJuyxlm5Os2xgSAaKnDJlkd10WBVAchZxxoJ2R7HUG/grPMJY7GbPPSrzJSanGy5BP6Jpz
LHndcMitjZE24WpJdG4GHTlsJ2T8DLgWwsIzYpDymCOPDDcLPQw0JzrmVH6wF07Rv8gogH129g+0
DVgC6f+/Z56E0qa+mXjJaAsKOkjOhGwQ6VlOhcNFIuIpZZl+GyWZQG8RiStG3ZC9bnT7/HzwUy0l
1Hu8DI+JqtAKyx84K51lXcFlPCZtxz+N8dzf7D8jezzEfR1tqESSYyUtxDd+7x4L16riAR7i72Og
H0RC4dwMY6pcd2jgiTmylEFfGSDvBmozCIEiEugWWj44eZmTej/hE1OAM0dUNDjfF9YbqgfGfSsD
TacPbRRoKvHSqG22JcmJMOG6tHHHwpNTCOqWKB8xxkfSFI4UWrP6p9RTy8N+ltMtkBHUufQdUY+h
H7o/3lNpx72Badkz1iUWLLtU47kYBKYTqixfMRZh0Z+DwknyBSrkW3UoO6FiaQerCm2P20rEFDCe
mzlv5AvIpE5eX7YzqUFVtF1D5ZrQiWYvU0xHlel0itvIACN2En2b9WQRDBuM5Ktm70MyeLemxR/M
TLgQ7JSZ6YI5il6qXQYhlThNOIXRcLnaNVrfeR200Z+mi99VDD0zZCDQKSkoYb7s4XoEcWvFKVzI
l1s4UrE6VAgdkyLnAcpH/EVZX++m5C5Zjv7kZn2Xr+RJLwa2OzFAoIIGhX88bPTjTGL+lZm6YsUC
D6cC3aLOdemFI1UVxbGFTYXQ+8x4domtKaZ73Iwgdme07HBdl/CoIKbY5j3XfGxH46xkm8HeqydL
+FIZ+dsnu7Y6WqiWvLoRTt2x0T5PHmbf9Q52dW/SG/WcOwiNvtS3b2PdtK98PjwjIUUq1+JkedNt
fY7Sugzz9J8pPoyhuFnRip7agqQbUXflv8xncMJBkNoh9xDquwgqYVaFwoPO5+Ka3KmTAit058VU
MVfQ7k5MTpSzKfqMHtQ/YEdYe6QXKRKfa272n6JqWBVmeBeE6jNh6A7jXK6jFbMj+x0IknYPVDMp
FXN+h71J7eouo0XwUG52B40jeFZ2hLGxiOFKkEiVzIMGximfxvLbHTlhSrZWje/75egHdK+RmlUY
S8ov1mDj3nhUlnrdQS+rE2UT4D22mYekMG1eZPvwiUnnCdbEDwUZKCUgX+bEz6zcEOwI31/wfi8W
vNpnPtLm84ke1bBrGEe0mBlAVEJbQ+8AFSwGSyQvRhk/9+etnb7z6VvZB6GtTnjzWqEMLLY91c/C
g+nlQvfbAqPn67SHN4UTAPzLbjnbzX9+paWEWpqPtvG6Si9IP2sBFcGVjybsQRTTcz4xCzkwYGGV
KfWHCWYwrFTj6M9/Mkr1xkoKWle2C12tfSM4eS+dENDOMNlNtcoBBfhfYAyNDgcXQTY6jeMh+Qbs
YzWZsAnu2lwj9n7Fvj9U1M4EJEVD9U9ObE7MGBcQKLP9hmkz3xRH2CUlw2ramiuoX3qopLS17I0p
Ql65gWh1y5WK8K/qOWdDwEXsFipqEiznZRrFuRqUF34tv8ofzpsfrZYILEc7d3NTe5GpTGUPTADv
t7RK/csNhCtE7Qdog4j7ahFXtTDimfcT05Ews439PGVDAkIcfZWNgNVi4U6+hEioOZNHOIxYACWw
Ytcfue2J/QLA3rsyUCLXMoRyOez2bGKeJd+IWQh2FBPhAM2a58iq01FbPTzffwgJZ8QbgSQOODmM
qnLt0vxFKwRKY+PTAfY5esd3iAqKJ1mvN+hN1TG1PCST5TD7/oeOV0+Oz7Y=
`protect end_protected
