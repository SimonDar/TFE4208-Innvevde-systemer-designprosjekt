��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j0y�ߞ��'DmP"l�8Ws����3#�P����P�ɻ��v�B�*����ހٗ��l�I�$JE�����X�(�>���'v���)U:���si����mY��������f}���/ p�2P�W���v�R�9d��$h�E�o���kI���c�z%�y��	E<|���Ur��~����M��`(���)dDP�>��B� G����Y���uj�%u�FgM4eaqP�}��=n��>�B��g+��v�a�D I�����r#�t(gò�*ow�KF��R�Ѷ+�9��õ:�K1�6ѕ��#���|q�ӻ*u,*��Pj��,��F�u����<�?�����C��T�P�"I�5�&�P4����:�[���4�dcH(�*��'u���}1E����(ʜ��)��@����ԅ�p����;���KOGl�~.Vn��e���NC6~���q��ÀL�{�T��1פ�s[Z� ��o���\d�c�DV�O�1���)��(�|�lJ��{naM4U�옄 ���4�k܄������V'�c�Q�r�cH�o0����_�$(�5}R�[P��RA�rIð |"\<��n�"Ͼ,{`qޒ��F甝2�h�"#
o����_Ĝ0
�#T�D�چ�㉾ڔ�0��o��)��!��a-�׵-d꒤V�(��ŸX@��`Cd��Aq�Y�ؙ�od1 S����E� X���{�ٙjK�O��N�s�6�R"�R���a@��]Ga2�'6�I��NB�Ǯ9u6Hj���
�l�6�����ӵ9��W��kʠ �2��6{��[FU-�p����"Z6)Y���6�7��T����t����5��V�(��y������{�ݟ�/J:���j��&Z(6t��˹����Xz�1���6F7�3X�.�H@z|u�o>�%�{~EVZ,f�xT�	yU�<�A�vM�E��f�u+�����_?�"��Lp�5n�Dƕ��E���ٴ�Dύ�X�p!I�^Z}���
X#?L��s�-.e�}�D�)��n��e�6D��<�M���E܁_ �$���mj���~n[�a]���,�b\���@�!ץߤ�"ߥ���&�l�
���Cv�A3a/@�&cꆞ3��Q�{�V�h�YP�;�dՃ\;��mݯ �;Qm֏7V����I�l�P�n�Y�w��ң�pV�"�4�77�[8����d���dU��%���NH��}^Ԋ�aD��"v"s�ӵ�6�{���6���۹�cu��P΃#��MHnt�詩�bSgl�Ͷ��Ɖ�a
:��5m��U5,p��9�`���+�������җ\#�r�1K)Ê=� �|X���C[C��o��3{����"����h�`�/�����sPCF)��yoY��x@C�" �Ud��#D�]!�ɍ������:g�]�n.�Mr��c�-��>�>��3&+@�1��b�c�-���`J�_�;D3q��E����@n� �c-F�dKo��^sٞ�ŕH|2B��dG!dЩK�w��)Q�RKr��!.R�1��֓Q9��4�$#��Y*M�0��������� wh�ހX����HG���l�Q��k]���;~mo�g�K������S�)�TB4��
�k=���qK�����4y�8P��_A<���/��j�9K b�&�����X�$���y��^�vy�%��v�A������<8��Q,�^ާ��H'<��G��9 I�;1�	 ���?Z�eq1ɽ�����d;)ޖ�n:]4�=�� ������޾����#j����k�̈́�M��f�� ��&f���c���K���R�x�w�S�n��'�_�L�<�tZ����(~��u�'{.*��д9N�����K^��`g8*4����7����D�#ô㿟�� (�~IC(�����u�P�����s�*Fy��'�����Qaã�䠓���K�o��E�,AIFi��{hr�����[v����Ϸ�ê�� � ROa�
t�)4ed��C�Q�j��Gj�1�{a
�S�`���κg�^{��N+��BiԋL�ɑ�K��]50̒���%I�"X�����nM�gd��SZG�U!��j�8��Wru� N��5��R�����o���.̅���o��E�,2VN�KY�P�|y<�XK�}B����l�����g�Jj/�`�2.jK|��z+��hȒ�O#�F/�����w,�p�����pdm�Y��w. [r$��~P�L�>� ��~�(WB|q��x��#�,��L�g��7��,�3x.c��qS͑����>z%�*M�I¦_z�p��J��"^���,�wl�"|�'.S!�NM�U��b������7�!����_�@�s� �M���챞'�l��^�v`�/�UuOg�H�G�7�V�q�J���@O�|<E�������:�ן�y#~j&��=��-���9�|���q�m\VJ�m��v,,8b����Z��
��c%l�+;+�(���{������O��:��f����:����|��Q������:8����k�Iw1Jt����Jt�I����KuhYAm%���@d|f!��oK����$|���T[u����p��dj���IH�Z0��L����m^봹ז�=��6�c	E�|bIjd������$��r�@U�Ѥr-�� x�x��@�y���Y.3r�=�k��/��!� M��u~V�E}-$�%�>:�:�GI���BN���kgK��M�ļ6�.��e�:ޘU�3��vB�ں̮K�Y�<X����6�\Ⱥx�[Et ����Ǌ�a�������s_tUƒ��а4�V���}�)�����vU��L�����5fwuP�� �3I �ivC'9�6��j�k����j�4��/Q٪O����rpqMX�+[��Ow���~���FM�@8#>����>������bͼj۶�{d#�YJ��LݷB!�Z=;�r�0)�&�XyGQH����rl�ֵ/����2���ǩWK�BU�z&�:�P9Άy�� ���</�9�����7S�)3@�B�2}��� Ӕ����F�#[�&��Bd�e��������6#+!X�K�ʧ	�(��DH�`��7�������y%���)���g�MG$�ld$Yv^�ֲn�A.��e������I��E�gb��PE��Ɓ	nR���n�\����a����H�;�X)�AY�_f�g	�gF�j��A���j��o��.��)�{��(�8�46�bd|���t�H��L���������c���Ёs}��"�-�ˋ?��o��U���'3ٞ�1����aSGц?Rk���TZ��"��8cS�_8��!��^���2�+%~y�� Q9��<�S�(jO�,� ������q�$�&l��ϗ��G_r�L�PJ.�֞/��ޑjiA��e1��a��CԴ+H����~�"���$.1<Z6�C��ؠ����"e��@��ʛ(��(o�9��g[��P�+�����7!��]Z�ҫ)6NY�\{ŉ�,�*�����]�����p��q5��p��e��=jȧّG�G�6uyp{��G�_zQ���M�C�F˪YOhj_9:9Bfp�ψ�LOm���@8���ǹ�x�rm��\w_2����R����h�1
XDu�8���l��)W�FF�������,�U����0�^���)w��l5�NM�]9�M�`V� .�Y���
>Z�֓j�%ukj�Л��u���B�?cg�m �B�@��d�ʜ�=�?jw�;����"��367����n�p�q*A��_���떞���,ק�ܓ�ev;q��<��+z� ����Z����042��t2�Xm�x����GB�S��P:�c��WG���������)�Ҝ#���#���
>���u���/v�������u��q����ʽ��]B�-bGԣ>�LyȖC��˓6���;`%q����Y����!M:"h5�iǳ7���R��a��Y����((���߿���k�b])h�$R�oл�C���w���߸�W��4i�x���x��������T�lvu3ٸ�?��Lث14ۣ�L��3�e"o�|G�
ۿ,��9[�8b�P�����߬�!�n��R��`c��Z
(+aQ&l��=��ޢ�=8�����<��)�n����\k/2,o���u��<d����7��*��Id�͹/��vY����9�;n鮥�̎}��S+�p+���>	uTz	�	���2�&-�rk*�n�$ G�k��͑z���Jm�[4��O+?�Kw����G�����ry�-3ѹ��q:��ʶt=�)2�7+��v�g�E�A�ꤛ1N�W�%%B�5�`5'\s���;��Y��˕MԤ��3�� ���T]��Vv�ފ@��K����0 DlAH%�\�
���
�������v=8�� o5t~��VV>'\�?�X��R<*
%Ҋgc���	 n��MY�j,^�t��9�v�Q���Z}T������i$�a@���x���𚚏� Wwϡ����e��]m������&硌�3�x�؉4����}8���>�5���U���\lĴ�BM��*���F�jY�7��+$j�)���i�ٴQk�i�.�<��������:If�;w��G���+|��]���[�H]�"�%rX͑�'Yjp��a �p;����<�wE*m'����hS$��$�lz��+�<]4�����++L�F}`���x-��C������(h�B=ǛmĊM�[��w���+M�Mil˾�$EW�G5}r)b��&�1����T�88i��K��szp�-4b��l�8uQ��Б�5���-o���}���k�>�Eb�S�7���J��Z�/�oL6H�G��Y�Შw�-�V6�CoM:_��ө�K
�v��#]OP������q�M�����Ld����znv��f�*'Y!�v$#͹	�l���z�t��qX���;���o�D (d��.W���4�U�>��mD���/X���W4�5l	p�����d��Ư��.q��&�@����\�M_)�;g��	!��π�~����F���t^ʡ���/�^��{mG���iT_��"J��R8jm��`�ہ�����aX��'+�%���2�!E R
�FW3q
����Y��iuB����Wn���W��O��{/����O�j��\qf�d��������r�GU��(�����kk��r�8� ��:Тi���I�G��V��įO�ncn�,t�d�밉
�Ĩ����L��|��a����0��f~������@4<kg+ʣ��C��pq{���*���d:��H����[���S���c�b�蝕%�x����P���t8��� �0�O䒮d�(�.�5e%k��v�\ �.$����˯�����o0+���]���Ӕw�2�p��?�5�ז�L�T�jp���k�7����Q��,�g��1��� �9�1d I砩�,��~��\�>F���ĳ�}`SO'sŕH�x����rn �����٪l^&��;ʻ�{��kr�u}ͥ����6������������R5���x$�vtb	����w�`�_KaA	!6$�$$�'���7/+9}�A0��*����i��]Wp 'Z��N���5��?�]�g����3��VЍP8kO��P�3V��4��p�ah�ښ.�Tt�CC6B�0��?�.�5}�SЧ��͜��E��@���!CQA�2
<��<[��d����C��@�0��վN0N�qާ�<�(0V�·��!�c��R�yǙ�;-�����K\�ץA>1
����c��?U<�=G��&_<��kT�/�Q9���{�*��G�`P9�n�)�\7M�q�����$ �$��IV���_��h`le�:������pp��=曇K�C&��5�\�H3��P����r���'�!n#PR#�X�c���0�k)��a;~i�q|���5z\ɕ`��?:N`h�D��ɛ�Bc���!G81�JT4��o�ɔ7�H�.���C��0�!������UO޻nr��=>+�eDʢ@��J`4���,�&�h���\���L�"�tu�'����M���q�@2�/u��.�TR��l*L� �2<��pڧ�<�`�>p���0�����*4~We��$���-�G�)\�+B�X�D��.9�h�Ų���P���Ry]�