��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~	U�_K�-����(�谝�of00�,�#ʵ�r�d���(��Ҙ�[�Ъ��ԯ�JIr�*��^��Lq��q�	 #ב�D>�gZTHiꣻ!'0hdU��*?l��B�Ei����Mw��D͇���4��|��HjߐE��C4�*�M��p�^U7S��.�tz%��wQ�c ��)����XQ���?y��_y��k�����}��y-rN%�K�~
�ţא')�� �.@��v]*�.S���3{�}�a�Bc|�A�%c@��"F�������5��ԨL��H�b�QC��S�`���t��"������l��,QH:��8����
�Cd��D�@N��+���
�����V��q��l0߸*���e�6t�)���C�����3U��c���'Q�S��l�b\���=j������Y�/ܹ�9ZYq`x�]mM 8��ANO�L� �RHAUW�e_O$'��L��
�?�9t���S_�RE�6�{��Pe[�˦�o0�Ch#�u:��;rs��lS�W����h�A䳀Ly�7��/nB^<����Nчܽw����C����s�������2s[H�!Kr�2�C��=���X�t���o9�k�\D�BIVϻ	ږ��Q�����H�s��ط"�rpN�plZ����Yi�H$ϭ6_�^h9��3��:x��_�U���-�T>���z�|��B,=~�cZ��S��uJ���u�B���m���J����m�&?v&z��B��fNy� ���k:F9^��-��`#�u:B�Wd�{�6K�#��i8`v�s&�;!L.��Ֆo�xf�-�j�E�=q����2��{Rָ�u���yZ�n4��,�$�a�	7�b��|:�I1�J(�G&]d�puji�`��L��@b~��
��d�_������W5��u4�v�AT���N��Oq+��}˔uB�0,,���
X/��Dafˍ� ����,��Pڳ��T!�(~V3���Bx�����B��/��s�a��3M�F��o����+Җ��t��
ҷJXZ���#�����s����-})o0+&���z]�u���6��n�,+Ʋ�E&��0���� ������ĆT:i�Jʬ!m��X`7�Je{�b�;�a��39q�G��~~�����#��s�j̒uq��S�=I3 �-���Ԟ�
nP�k�.��M�u�gT6P��!�С�M�� �F��CV{��L���.�vJ����g�P��Ƿ5�ynu�U���B)�`���Y�R=�647(%�D�f�RKf�MI���X�?Ye��.��V*��<�̻��5�$T�cs��U�Љ���Q�N�B$��,%|x<��Q(.P����8�=�Lc�7n&���$�Q�� ǖx�O2W]i7(��☦�$��k��TRo����0����q4�?��)�h�§�\�Vb�F��B� L���%,z%S-������Z�3�e�u
B�ۺޤn�v�Нxc�i��c���}w�$�x6���_D�w5�x��%�̀x���u�P�Dq��D�@M��4/�W�XO�%z,
sb\-�|���U3=#��!PA��XǇ�[[Y����3ƣ�~%���CQ����u!����r���>��׷2x�a���w��gA��i^"r��ܫ}��`I"F,�y��*q)ln�§Fp�1O��4��?���~�,��R��������
�|蟐D�m���{w�25�*٬YP���(�-%B�Դ��	�B�9�u��������΅�Q �]�����RL��e�mh��flY:�E
�68��/�X*��pHH�y�J\?S��E"Z�{Oж{,,������8�d�-�	rU������ȃ>����C����`UG_�e�"��P��i�ןz���C���c���`m`D M�� DH�["���҈���
�Nn����cV�CՔ�@�=1b�Fa���f�z�40�K� 1��ȸ@'�.�Vg�NL����.��VH<�`F���&,m��u9!��gR���,Xm���v���'"�sd5�4��?�鉙���ΉS����4��ZOLC��䦡���*.%˝ݝCr�w�4?�GĄA2d#q��-�v�!e��|��i�����3,���v]3�>׋�Nj5����QG�Э�p�,�	��/����pt�8M ?��v�{P��0:��	e��1�-c1^������NJJo�4���$�d�k��eI����O ���y�/"�E��3R�I��M(��|�X�I��}o���h�0�^�'���'8�0AF#��l������=��r6�"�~)�����h5�?�>�q ��إĻ���.�%n�%�#�m��	�+U;I��t��5���T'�9 Y�Yd�Lm=$A'!y���Рc�wX�-am��
$�s�u�������m���*��
Q�D��yơo��jp�ܧ���:� ���2q�s�Bػ���"� �����1п���������2]�#t� �O?�c��8{�A��»��%<71����s��ĸ���z�MW�(b��;M�I��-���n�fss\�0���m���:����ʓ��"�t�c"s�5�Hx�^�:;��4N��!��Uo*M�s�՚c�g1�t���P��󒼁7�����x�݄��~,��{���uE L|WMÁ�52@K�
aX�B��ϐ ��u���d&�F� �hz�D'�&Dvh���=q�J$��+_}�=���}���s�s�0YG!�3��ؓ4��/Li�"|/�g�	���A�ߍ��G�����D�JA�+^b�i�����Y�������}�$��Y!�'�%Uw�D����G��7B��1�@ �����y!$cw�~��q
PHe�A"W]�ιP��w���a�	�NT���:P��L �&Nϊ�cTJ����~�I=T�ܘ	�;��^���/��$G�)��F�=)=p�C Kh�j��#�x�4�>%����ʜy��ϔ� ��(ke���`E�Z9�� "2����v��#[Hu��LI�`ȽJ/z̶+<b����E�}f'YY������=Hu�"z����C���a�ׂL�k�������=o'\5M,?�s��G) .*����5UM���͚z^^o�յ��	�z���b=Č
E�+��5����	�1̖��e�PF�%��,5���N���3�W��Mo���*=�22��V��8��t�q��m�Wp�t?>yԠ�YHh��2]�_�uH��X����?o�Xz��m�!��!�s��9��Z*����b)a ��)�3�c�Y��}si"�_H���!���o��7N�p7�<����Μ�>���5h8˿1%:P��U�*�Ȑ/J�!��C �3jPq��`�r�w2&���Vӑ�!@��t5L�P��?��q�K8w��R�`ҹq�䗚V����ޯ"pz���Kc��@�,�ʺ��5Z_����-�v
�p�X߇��&d����_Wd��BO��AZ�h#����^��jP�������̑R���6�3Nm��v�Z�h�pF���{]��u6_�|� ��R;S�ҧO[�+ޗT�:BNetk���<㜒�3wU�K�g�]�*�i�T@^��О�B�+"��<��f�k�1�^�s�e�K�4����]X�ʇ��vم�w�?��U�.��
V���Hi.o�#W%^y<����ٌ;�|č;C�eץ�К��oؽ�ؤ�i��?�QG��y"`L�6�)�ͪ��N�0�ތz��^5�1�'���ǸE��Ûo� P�^��c;&�����*M2�|��hUN�J����K�ҟ��z�Ӧ��W3T��Ә�� ��.)�>�z��.p� lU/.���F�ʛ�h�t�R��D�4����#�{�!�u�a��
��XFl�͊�4�-3�t.{"Ț�b���.��*o1��	�St?Nڒ�',��>38Ǿ����բ%A���l���!)*��H�z�Y]�=�CC�ƽ���+��5"�����C�+�f7���P�Z-�2��27�;�0�~"户�,�0:�k�����H�L�bl9���%y��)rfq��� �"�����!�x��思౳��6C�)AD�?���]��O|#ɔ9p���d=MW_�[�ŪV&��ÿ��
��_Bض�I��q&�R8�|���]��.�Ђ�h1eX ̯�9T�_��_�6�g��ؾI��9�YK�0�Н}Y�w��p��f��#bph奇��:��f��P��X"��WARv��Z�W��{?��L�Άw��q'��nE�h�^��F�`��1�0H�	���2<���= I�^��R��A[��Y�V3ua�Q�nE�-�C���#|��%��+�:1�9�R��)���͆ˉ�J�:�Ԁ�V���e��l+` �i�\�tNS��IG�M,�]箁QȪVt�3]�7}��d~ ��L�ߘ߄���&Q�p�e��̤r�#�,���Z�W� ��X�q��(b��`�%�r:2?o#��vX�������-p�mΣ4�r��v�t��*pt��M�a�f$׃b��~A�p� �tD��sFB���#
�����q���c���`2U�Ԇ����cی󋭱t�Q����^-����{6�;GCn�@2"����b�O7���]jNgW���������ʑǈ(|��!�#`��h���<#kG��"�{�5O[�oL�ߪ ��k�$f��"#����4�V��bP�m%��s�E�T.�d-@�\_��;�<	��!�<�4�"]϶��WO8�܅��d�(���}��!��6B]4�D9�n��k�M���$�r�+(C�u�eT�X���6^{����(��5]WK|�`<���Ȅ��Oö��ik]�D�_���1�B���P��E�!���&�@��F�O�l�vo1�1��0�O�w�&�"E�!G��,tӍ'ɘ_߲�[t�j:(�F"�+����t�h�_j�D��=<NN�,��
�xq��d��I�U�?��w�����z����$�4U#�)�A\{���"�G ]&�6j<�4�{^�B�=�:�K�����K�OÓ�Y`�E�\ϳ^�n/�#�հLSLd]&@�eM����$��ӰV#���x��rʶ{���^f�Q���_Z F�C	�i�R]�?Ƚ�5�|���H75��A����k�ˌs$bJwx��L���