��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U@W~z,r#�9˨�κ�B���Ԩ��^&����ם���/�8ai�j<�@�p���m{"��ƴ4��w�å Pw�JM�}�i�Ƈ����Jf��/0$�}�C�S�2���R:V�������d�61�חy�N����[V����9F��� �(��uixl��q��l�N�
��|A���~��t�e^�,�I�qt�!�]2�c��~�c����#�ýgf�jP�]3fෘ�/f��ԋ���~d�r��#�@s]5�A�=�b��Ҡ��v�icش!�	ꏭ��zz��� bl�����z�)�B6��kN��Nc/�$'��@�S��Rb����@GF�(]��AzW�"�V�I�E��4�&�p�Y����k�M2�fe��R�!�ןny3x�;��+vA&4��|,#v�R�(`[��{�� �m�os�b&mH�\��:"�oх�
��e���a�����娥�`2q�*8	Smk�@�&�#�G����ws���D������t}���	�ATuf/�ʸ���Q?��(\� !j2ҙ�1�`��[CM�X_{ $���:�ٞ�A��lj�7�d4�?ItC�rL��^n)�7H8P_��oEf�c{Ɲ�$��Z��:Wq����{
�/2
s�))�R�J޲���>(2h�L� �[����URE�ZS{�LR��Qj����ZXn��S=��$�u��u��<������F��Y�����Go�H�����PJ%a5~B4܂v�}+fٷ �xϲ*������^�(��)�Q�Q�EBa���y�:�,3Q}^.Z�O�jQeYX�>�2�T0�/�ʓs}i��e�}�nA��J����H\�����ŒE�~6mp*bΏ0 <G�4uJ)�T����-q���ܥr&VY��~@ZZ�:Q���i�o�t�"7:�&�
��Zh���� �S�G�ZǞ9�o�
����f6�Қ�lȵ�V;4�60�89���)�_
.ɫ-C�(����FL��*����ڡC�4���Pرƞ���(��nn���ALN�&9,-�O���9��EO�	k��bؒ��eȔ�ċ�zy7�~��z�)7d��%�^7��R	����>���%�$]J��H,7�6��9�c������}�>3�w�5��v �s���Lm0s�D%��ӼY@�!GV�&���KB�SӸo�M ����c��df{K�T�#B�>�ד�(���սFa�Ѭ�Bs|I�����h^䄭������4����,�=�ׅG��M�+������dRn�,5\�#,%;�8��;,C^M��Wt7$7� Q�[�Y:�D6�cݴ�h�)I��U�r(^aUfq��t���!S��34f�J[)�lh�����R�82O�ުV�<���~�}�Y�w[�+:��]�<qD���Wy8��D�R���wI���@(DG[7�8�VP~��rS5�,�IgxьM�Gp����㊵`>�5��x嶽�ٝ]��-�) �~�/�T�Đ�oBs�f��J�S������I��'3o��]��X�>���6לǖ���G�ϳ�- �>OS��4YYD��TJ��޷�P�x�m�;1�[����FX��ᡧwGw1��m�$+�y�C�B����oS��u�����^�������s���I�L�R�-}�fgN��oݣZY@��Y0�l��s�$H�.���UbXF�T�ǻ��:QL�| I>Չa��'Z���1��|��N��|U2��dlEY�]���s�Y�k��W��g���4��� ���Y�����q�2���Q�Jzsl�� ��EM�m\an�z߿&j]�j�f��wy'���% *��g��}}*X����Ǐ\��Ҏ Hhl��0�O�}�Tw�w�+Y��~I���h�`�����W)�p:�o-�i�y۰���԰�f�6��ze�5������a��'�ƶ���g��XY��o���U>���� ��.��1�}U�L����� ��!�)��n��pM*:�q�s�������ZT�B]���!@�!�Y�?e����������9�ջ�2��9)���c�ܶ�Y���N�;��<��K�z�h^�?����]��
~S��G������qƌ2��誰@�
���1��o��R�\vh��%d[`얓ǎ;.7ƕ�����Aalb�Z�����Uʰ�r�Md$�	G��[䈔R����.�n-�[�����MA0Ǯl"�n��up�c�C�4���	Z�?5�E�����VwP�CNu���j6U:z��C��_���B���>�}on���U��C���5�!Tt�g���g�3o��):��u&�|�s��ۨ<��]9/�;wե��E�΁��=a'�]'~q�!��*b����^�V�����0=�?�l��D���s�U}v��3n[�q���]�I�F��n^����.�
�A�T���hኯ�Yo�c-NF��nu���ዠcF�wwZ�Ba�1��x��}1ώ �i�N�X���5���U��`�eYc��a��H'7�N��pt-�c1���d��:���=IuZ)8�$X����oBX=;/r��j7�ְ�y���@�͛�*I� v���,Wi�iv5�SR̐�N��#���>�q8�a/u�tl�ߎ҂h*(�7*i��(����rk���/�h��poӢ�(\xM�
���tT��ڨ�/f���1đvzM�^UI�����2s��9;��}l���Yd���x�7Zr��.�H�	޸��~��cƭ����'��Pm(�/Gy�5W�M�=����N���O��i�t��Ⱥ��$ya�C/�D��]�26[¤�nL��Fn���gu���S���Z#�GI��tH���J��bZ���x�;BkR=b0���U�/2�?^���:��[�m�4-~�V���h�V��S*1�E��]�$�}Y�nݥx�O�r��5���v�i�J�o��o�ʛt�k�~=��ͼU��O�� �2?=�;��6Cr�f��ZRT[#^��b��=�^ޤS��~v�\(m��+�$=쐐��m��,v�'�B�E����m\�Z�o눡}4���+j��w5 3�PoD#��弜6��`7f̐:z��S�����0�=�T��r̮&;Jj�Q��I��uf�R�[EE"���b���&B��W
D؅��A=�����V�����	ܫ��}5��P�f��_5����¶M��{D!�~��o�K#J��1��^u�ڬʁ}��ыjH��Cjy�0�an�{U�q���@��U^���3� �Y�d����H�h�r���w��Dn2��p/[F�������Ny�Ԍ�D[b#=���R��n�L��Hf7��Zb._��W�)�[{d�[��G�7�"��%;;=�]kb[�;+Bɡ�q�z��3��*9$�Y���P�-�!c��������,�Z�;���yv[tz�����)|jZ`i�YX���5�f���L`R�ܵ�C5���QD����l	{j=�S�?n���;+�8N�F d<�\y��K�(�dO�)m`�ʢ�޼���.C�������k�iI��+�;���ca
F��zN�,��1��|�������{�֓�\MK,�O}��P��X4����5%�t�7����x4�j�Q����<��wN:D�Y|}���^�-���_�ZB|(�˼7~���*
� ��>�j���E�Y)赵!��#��e[I�k[��ǔ�l�� i���/�ar�ʫ�9��ȵ�m �(�IcI�@b���u,"��vKx�����������w|-���b��lú�,K8�r1���ʲ;-�aG�j�|�̄���w�*��$_0�%Af�'���oGg��\�sNKK�W)�	ST��]?]g��aȦ|6ύϮ��wm����xB"=���D���o�/�fL�q���;�M�:��*etJz'Ӂ2?5é,����g�&|RS{�t��g����w��;�?o�VBV��p1^�� Ŏ����Q��s8���SU|S1�o���I�S�W���]H���o[!�|W1Q��A[=�����"�����&kKxs�M»�1޽��i�?f��	=2�`�q��c_c.(�����r;S��R{%��=a���ߺ�C�Հ����w��1���cg2��ܴ�b�F�}��z���0��_H�W{�*� 5Ѭ��]C&�t6l���(Jeo�:�����` �Pd	�6����L,��#�K ��J o�J�h@A�)]��֮c�L5$�:�9ȽDĜ�Vm ��B��e�S�JW���yo'�W|IuG�:Z&�%�����ব�O����:���4鞚�-�L�����,KŌo����������7nq1�K �t��_^��
>s�'S%��/���13r5�zWw��JΖO cf-]?9l�8��,��O��Jx����
^&N�I�}�}8�z�/!Ddz�#�VR�IQ!����y4��s�*I��)H���G�����4?�F��g6�Bs�`�8�`
q���)�f�x]7$)��BZ�U��Ev�
ɡ�xĔ}ů7��tc|fK=�0�<~�.�C�E'1�	Ⱦρ#���U�Ie?�
�r�T�hu)�?rO�G2����"�OV+c#�Ѵ�K���aDt��,�X�\��u*9����K:�F�#���7��(��2bm���jj��g��a�T��:g�v��ʹ��&Ҙk1�+��qg�A���Q5��W
ujK͞>�.�H�6�D��n/b��kD�n٢b�����|����'E��P.hT�����y@�Vs(��D�u�:�a�|�#;%%Ȗ���A�s��5����H��M�?MЭ+|8��7�*nhWCRQ���yb�lA��AE �U�Y(U��OA͑���r�_�>�$��s �Y�˾��OX��~�JHj��g��@����ːH�4U�T\��<��G�(�q�S�桋C��+���X8�M&pM�8��� A��jCL�N+)M>��,�[JhPe�mU�9�|o�b*-��S�4��x̕�.ق���3�����C���p�H���Jy�TtF��Vר��qw��1�
7�Q�Q؁��2gU�WPU�
��Z���,�t�T��_���%�_�#�c�I2v{��Ȫ��J���dd ]�T�gŨ�F�<;��_!��+'j$f>�s�a~Ҍ�C7P��I�6J��KL��'c�t�Q��̣��R4I��NaT4�nMh��iw{�֊0e ���K!V4s�9�GF���J2t5iO��_T�1S��ڿD���J�t�>x��n�x�d1�ޜ�|
�*��W}|�hڀU�..�; #���~�1��9fN�>|���P�-��������g���/f��ۇ5v��^}л����U��<���w��n����Pm�bJ#Z��7�m;+�y9'g�l��K���)� ���+4�w|�Mxh��l�|fxl���kȯ�"�5i�B�of�wj�r���TG��˴B�ZƷD	=Э)Q\&����sPy�.���7��;u�L
��>ڈ��+	�̖j�!����^�S9��֓i�z��E�"9������qw��6Y`��k��,sZ\���x�3����)�b�j��Z�-IAQZ��y=�Q�x�a k\�i��jZ)��׭��c�ű2ǝ?(QS��]��XE�  ?���1t��g&��ߙ�t�X�]��;��m��(�61����4鞞���èGt�I�o���7G6Ko�!��	���}�hc8Ela��f%qu��PMԫ�~6Z(���O��n?�m���l��$�'�DP9fM�4X���0��挍VK����^n=��\2�\T�3�;K��n=�[����&�$wAl4i
�T�'��H�($Ҝ(`,�,_Y��{�nAm?j(����@������B/*���EY�w�g���I�uu��0{�z�7���EP�F����S���H폹�=$�I�1SB�>$O���6Mv䌌�ܢ���Oړ���_��C��C8��5�;���̳�=�AK��U��Ѥ�9"d�ƺIvnH9x�3�(�{��W���á����Uv~W9�}<�@Ɩ�C�]�)�����T�'j��rC�����B8���n{Ԅ���KDG������<F���?��}�R$	�����W.u��zM�Uwǅ]!
vf<�%{y�(D�ʥ%6[��������9j0��^������Ib�b�إȈ�����S�z���t�n���K�#T��7v�&�\J�U�)�1�j���Y�'����cQ���i����\��h��^��nH���֗�.�J#f�L�0cY����:��\���Z�d�t~���{�T.*�`����H4??n�d���o�e�ib\X�jL�>����h���7�Y�X:b�x��<X��1ll�C-
&���iJ���r�ͫY���Uap���1��j��9�vd)�G��3���q�=d�#}m��� d_�3�"dK��x'##��C
�s& F�����f��0�c��'F�8��2�C77�bd��@���9�*����W��:0���H[��?����)d����M�u%�]͗N;&�������w�R���M�@D���t*:S�q��ea/�)�Q��/��B��V�j6{w�[[�V��AnNչ�F�a�)!�ܩ�9/1�̂�ˊ��3椾�YgG�o�?�'Y�{�]�E\Q�Y˯v�(��9�?V6I���G�=�%@ĸ��W��ۏn'l�@����S�k�.ޟp5��u� �6���4F��ȚK���t� &�Q��QrϽ��ܦ�}*�9I!驩eL�ֳԾ,O��q�[͜s�g5�?�u�F%�/�Qd����1�%��\.�˸6E(K�r��(0���0�#Qw���$��uɐQN�	>��N���u���\���/�e�Zz[��$�����I�[e��F�h��W�%�>`4z��nF���)[.���ag�Um(K^,'��jmZ���ZČ���zU%_��7�>
i3ۖ sCђ�����14WT�5�����m;lvwY��fG}��?#���dT�H~�es��5�.1��V�q������;�%t}7|�7�����ի5��l���_)K��[����8�1�4�By�Z��d Ϧ��ԕ��Ӣ�uj�=�\����a!�����k�G~/
����-�r�/�D�_��X�8�ِ�B�Bۅ3\�U�Y'���>��~h1�)O���>�I\��QӮ��t�
��T�e{���L~K���+=0��DRN�'3A{��@N�<�#qTZ�c��(�сkCi��3�ɟWI��X4A��0B�~T�
�6�{�ހчl|oY�aqiQp�\؅u^2�}��v=N��d��V��ߟv#�i0�i?0CQ�S6��!�Ѣ��jƠr�$H	8+��a����$y_���T��HE��I{��Dsְ�/��/��O�Z���o��]"7��H��7��p\��SI$1���ěz�0�+��?Pi9�=fvd��r�Ё��1���L0����r����o�ZO)\`G��qi&0��C�@��03��|�n5�<r����0���<��q���.%�ŰMo\�𔘖�Dz���(sq��+��&�3I��W�d�g ����GM h���}F:䒷,t. |����qq�AK��i#Ql(P��lxk%�4zo�NW��~y�BJ����ZB���.���Urk���~�	�"��N�*�i�z��U�-iƣ����Z(v��ʣB�?ɼcYa����O����3�������:�P֬��1-������-I��vR޸
W
���_�Yu�L��Ħ����E�׎NO�ݽ5��� 	��M�����S�� ;�H�/2s�^ͦ�[�� �01��got��`���܂S�@z!��ojo>��ϊ��cf����/��	���+���(R_�z��[���Mr��"�G�1"ݖ����x0�i�-3�����F�����'�lF�D��`�9�f+�t�S��{��蜛�.�J�������6������A����-��J{즿����73�]�>0����Q����D^�vP ދ��S+���M�A!�Җ��+X�e��� ��H��R��o�F�WL+�����qzR�U�'���Q���\ZQ��ڔj�H�:<,�G�f����%�����^ɾ�w��b��/�l�0Éo{ <�z�緅|�ܘ�YF0�E�7�1K-�3�!���� ��Z����&����]�޿���0xT7"M����=xĝ��"H�+�K���i0 #���}*,/Ѩ��0(��;�?�6C�u��\}��ۻI���Q���&�`���|b��2��4����w����)�kQ���݌�:�ν�HQη��}�@��P�.B��[�p×��{<����� �
��s%3�Z�q�o�T=�mF<���w�{�m��v\b�}�U��Z ��%����4��J��ߦ���Vl�ExC�%���q*1�ن99vDX��i��zY��`*��Ľr���3�7*l�^��5~k!Y��a5�tW#�0�(�;����[T�1
��i=z���A��MH�� -�i�Ґގ�f~kH|�fH�m�H{�a�@|�� wЂA�R�D���t�r�~�c�f��OM���o��q�*E|W�e��Yq3q�@JBl�VX�o�ps��(y:�k�G���l�	F���$=Y*��'���^�6�r�80�D�]��uĺ�b�!v�|~�P��X_�k�����M:;x��,�C���\�P�橻���X�l��F�,��Xj��gx�M��b3��R�a�������a2�-��^��ᰑ�	y�q���0k�A��;�Ըϋ.Vxz��8���s�zhօt���<�V?8C%�?-f��=��#C�-v"�-/4����}ļ����Lv2����Z\^&�8���*�wb-4�	� ���0�����a�#� �i�xE0G�N��I�a���=���j2W���a\TZ�n2t����;t0�����Sc5������f��ID΂�!��4V ��À�6�����U�ˌg>�p��5)e����Pѭ�H|��O��⼞I;�آ��uH?P�$8��UaG� �� k�A:��-zCC��x�����~����w�d&��m�H^�Dܥ�B�;9O�}38=����^�ڛT%Sw�k�(5����?��*m `iޔXfp�����i�u���1s�]����y�� <���!{�����61�?"�;��o�=�q=/�"���{GS�aK?� <P�{6�'0�~�j"�Wҭ�����ڝ�����OL8���"v2��:���	bG�A[��*�bw&���Uߨ�1W�E�^���P-a�� ��c��})�@]�W{6��N V�L�"�bYa��	zf&e�QC���I�S���_�^m������w���,·$�-(��Ѻ������c�w7hm��p��n)�t�����-1_�	'�r��0��{@�0�&v�a��}Y������1��_C{���*���ﳏ�u:K(�!{�	1
<V��J������Q]�\т^��n�6��W�[:�����	L˿&J߯�df�C��t��.����~	��]6+����0rW൯^Ii��p.�z�~��~\���R�}`]�����ϡa�}`��Z_gM�ŝվ6w�M�R4�C��iYRp�q�{[�|[������~�wf})�.���a���(�i��*��j����bF��0wҮ����ۺ���π����m�i���=���Y=����F����{��F9xt�8��^Z��j�Y-�Ut�l<15�����F���<.�c	ȷ�զ�����P�����%�{$G1�\ZG��?i����[��N�pM�ߺ+�\����]z��R��Rf�}M"�ͅO�eIM��0�{VNK��Ɯ�©%%�M9R��L�	�y���W�Փ�+�����=0�?�ws��ff����^�/M�=�� ��5?��>��-�I/��#�ԗ�C����z�b���U�ױ��(yĝ�ط��'��6�E����O H��`�����f�l�RȨ}R�kX��}z�K	���G#��l��Φq|b��,�\�Cg:��$�ɏ�J=pX���Hh�$�I��>����-�qh�e�����D-R�&3?�Ic�2s8��
io�	 a�H��
z��!?��E�nZ� sx��\�u��A�Ϧ#��T����{��n�ب3��J�O���U�%��u���&��8���N\�M?s��9d�2��nE�	�;/t��	0V�;=9m�2�'n��{l��� 4TI���6��j���i|�~�hf���C;@:���d9M$\�@�ϰo��V�VQ�Pd�OT#��m�;fT	U�˕��M�������4U�%��e��J�:)l.�oB�*	�.%rUp�d��Pq���vf��|�Hu���k�ne�����������`3=�J��D�kJ[�4���C�Ț��j��"��r'LG�a`�BG��9��Z"�y��Y��� �VY������{E�������B}�P(��	�ɭ���E�Ԓ�@뼛q
&�B�4�F�z�f��e�&�Փ����=~6�dنF�� ������Rwv)�ΧR� t:0E����ۢ_�n�g�w���P������}d�̜�����o9A���J�O뱝�̂,������%{�&&�~�p�'��;-�T��"/���`4�cb�[�än	4.]N���K�C[������w�$t́≄("�W ����U�D`��$:�"?�rM!�n�У���[;��?�.PC�0�-�8����
�Y�yj��z��H��@���g�k"F��dO���}�Q�>�� T>`�<䈙��u�E�w��-�`�|[h'q��nz��b��V���\N�D�R%
!�h��ůD=誤9)����}İ�24����)z>c470��>��6��������H/-yS�½8�����F�"Ct�	]Ǹ�e�
��8ijS4��:�9���[�.d��B�w+f���5�U��u���Qn���&��D�{�F�B,�K�6D���e)��xu5פD�ۙU�F>o�w�p�L+0w�^!㏨�W�ݻ?^Ή���n�ѓ���>�����qM�!7��Q-ʛ���|XK���~\�����6 �1��9w����eag� �]tx�C�A?T?� �g]iPko��i)-6�]�ʐ(H���ǻ����E��%zd(?���Au��Ȟs���ۄW�O��"J7ݩ�k��Ή0��)���T��%?8	�l?˽"���������x����G^��\�n�!�B m�����K��%yK�or�����bxQ
_���(��ܒan��e/�%��w�'}c_-�唒|�m�e��O=�nk"��9!�`"xu����Q:b�����,p�L?��j�:`�Li~z���O.
i�D��K�I�r�Jp���%&�}�{j��LA{�)pn�q�[��Hڤ�j����F�y�d߫�C#}@�^�U�S���WFFxt�J3'HiV���>�P�S6���-�*ȵ��I����ˊ8�|��{w���Óz��09�2A0a"1I�-����<��_����B=�t���<Z#紹�-3���${��M�M]�;��
?�?�yd^-nZV�s�@Q[���C9+^�gF�.[��̩φ?5����Y�a�¾�h��Z��<��⃊���X���j���.띡��v?K�XB��kl�R.�Ĭ���rS�Ӌ�4�0|٭��G!�H����ı(bQo�<�OG�x(C��7wX�1 ��;;�?�c��Ա�Y$�{��Z{��\��0G���;��lC��t����u[����c��0b.�þ��H�Wx�	Dہ�wE��>kK����2����,l�!>��uxY�x�>$�iVh�����餣d*�A��]��M�l�ߪ>�D�l�"���ꏛd��7�Hd
�Z��"���럕�ɡ9̄^�ًn��æ�s�ߚ���c��c׏�%��%�R�<g����va1�Eo�Q��]�#��gA
,ۇ��,x�ZԘvC�'d��|�� �u�S3Ď��}�zX���������nJ6��u���B$�g�ɂ��I��lRB)W�7'�xـ��͊zm�Q3�O�j����n=�{U$'t�^�R�2�@V���ݒT�����tiu�	��;��%��C`��t��`q.����C��+��:0��X�}��*V	h�[�{�������d�/j1�9c� ���:Z
d�z�J"�^`i	#�_6	���NЈӧ�o��1d5�(¦
��ꘐ���3��]�+O>�U�e'�hw,�rgκ$��uF�*���_z����Zt��u����~�T�E~���`גDR��g�=�4NPTUo0���[�<��VI�n&!Άc֦ڥ�=���m_��C����"���M�vT�	�FE栾���PY{�{���5\��iĺ���eZzGW)s���j�ގt�/���d��j=&��h�[M(�[c��}�b�ko�=�dnO�F�Х����@���m_}����.��neL�0[\e�7�mH��������M�!k&�<��J�SG��6}�ʧ����H��'�'5�?<4�W����V�&2W��YX����%��)���=s��RW2{�ƨ���i��,s�e�Ĕ��s~@��F�Rώ�Ǻ�����p�"M��N�Ȇ6x�d�pl�g�/<��"�𼀍F�g\�Zzb��V���P���q��4�Ԓ=���չJ�O���<u�(Ɯ�}����{��RW�hՕ42�b�|��=��ٵU���Dy���{	�s�BpW~�#��� i (�}����UA� ����ژ�y��
�T�RwFX�Ȓ=`����B��#��vF�cZ[�Y##�C3����J3T�L�.׽�
k���Y0e=HBA~�	+�i� F����l>X k� `
4��mR��鑍3�Z��¡ި�q�������Ղ�>��Q4\����E�E���b�@�T����w:A�#�l{�Fː�č��bT4���fk��;E�/�C2:�Gfn�c�/�x�zj�qMO*4s�<��̉u���j���Yo�#��!�/�yG �(��6�:�8�2Zx����3���1Uz${���_A>�q�;]|�F�\��u[��fE��(��s�^̨��D:Ɔ(���9�#?��4�,�#[�~<�߫F`��cĲ.\N#�S&���� ��e�Bf������
i�4�C�Bn�H�1,Km���mT��s��W9  !�:_��'| ���a�Z���p��I�(��,��c�oPxU39@��ѯʳD�#�rB店+�
�7�~e���=jP�i{փr03��V�s��<��EI�����玉���q]�eг���~ �>�b·��H��R�˂�Y������Y�p�����Y,�����eŪH���	����w��}��o�bsV~"[,����3^����N��*�!�6g�f�\լ�4�hr����{7�6 1��e�aB��S�~m��3��J�����N'��vA�k�G���RS�^}���
"�a4xa�i0�(���-&LyC�yоl&V��̊��<������|o[�N8�U�w0��}��Y��:Jm��֓Y:\�{��m���<��ӆO���Aͣ}�5�n?l>�PV�Ǭ���D�����_*���G�2��sRۑ����� ��V�U��FW�-PVR-#���O1��r��ֳj�����ԦЏiJ���������<�� �4�����2A p����������>F���髰�u�U�r��Γ�Q�A��Yؒ>В۴��aJ��¿ه}ǆ['�P��f����<Ǜ���ә�b��@5�����6]�����
�)/�2v�Q,ͣg�O��}�8��= |��6�����*�a�����b��n[S)��rƨ�i����\	�Vͼ�1��H�H����i�8��=���B����
x�n(���e ���j�9�J�Gdk[eO����bD�ht�i'F�������]`Ϯ[���F�u���Aq`V[��z�����k��)�$Ѽ��[��t�%
�L���l���
^�Ky?�2�U��#��Zsq�f�dr�p� ]�J��s���.�^^./�;[���i���|dG2�M�:����8�5�b3pl�7��b/s��8�Y.Y�ιUԪB�/<Շ�e��R�M�x53�f5�h�o!帏욯b��J��ǍJtK� oSj��/���e��&8r<DҐ�[��i�,�N�8�z�|�㙂CF+��aC8���-=�S�kxn�q0�*NƤ�%c!�`~/�yYC;�3p�x�(�n#�-K<؇Pg�*qP�u~sCO�o�5,'��2;Œ�p5S���������*�GR+��,�+4Ф��x�<kɰ(O�5�Q�*���p�LhMӪrU�:��^��gi��֨Z��l4�E��#�zg·�)Q�V	��[8�Z�>�sV��W����1�La��#�51n��-J~��ӝΪ#��yUu��«�O���I�ޑ����@;��WPoj�b$L�;���� (B��n ����YL�a�$����`U�A�jj澮l���ߤA#�+>�a�`�2$��j3�Z��]o��w�b�R��wu�%,�S) i2S9�QL�f�� �
��5��s��]�W�/�K[K�ʝ�z!�D斒ت�z`�2[_󣠐�J�)	�e�d�q$�����a�/�v���a��4S@j��A�?�����zλ@��#��� ġc'��#ej��o���Đ��O2 ��C`<$j�c<��n�Б�'�J�)���Zr	.6ݩ6�f�Y迦���tM@3��"��GkOgz�~��}������^ƃ����O_%?Up)K�k2A�~���������3����I���a{�1C�ea<`������Q�.��H2�	��$A ">����_c�͜����z3�fsi��4t�_�w-U~�����B9���Fc�M�$�������͛׮T��ifa�<�ʼ�z�~�(�	�JL*��${c;��ܝc�4�� ��K�f�|Qs�U�ǝ0��KV� �g :U� �+b�z�q�$ �۵NrE�0mJ��\��<��P`�'+��P�[��I���
e���j�x�X��g����v2��j�3s�|���j�}��[߉����oZ<f�����+cX�w��".����3>� o���|@�
{s�3gI��R���`)�)g2�5yF3Q��$?���)b�e�m`�/p�|��ҝ����P�4*�sHr���1˘���E�|@ 0.L�!&�g���I�^Ͻ�Zbs\��n��`��5o��d&(�b�'jZ�6|�Z/8T����.К�j����ލ��1:��9h}�-�3�pE�U�:��Xk!�f�)����;��vDDˊ�Z���e��bI�D��n��Ɵ��"��u8�)��	�2wp�ȸi@�	����3�ty����T�z�ە+L�D�K'����Fbzǐmo".X�e5�Iw���ϴ0�>���kȦWݐ)��e'=�2]N+ʲOV���F�[G,�m��W�T����z,���i�ї��H�m�u��j�]p�tc-0�f�p�BNɝ���=�Gpߕ��15d�
� �啤��>�f���R�O����vO�u������آ_S$��>E*�a$����� �-+�(���[��aD
�.Ja&�OF�Vo��<�Yn|�t����d�݃N�����=t*����Ep�#5���g�E���Յ-��U�������]��[�2�ܲ ��
�����B>�m�hTjOB�-%f��'����I2O��R����b�Ί����yw9id�6%�QH�]�?}ߕ:(V�v���r���i��ә�����V�����94�#Iw�J�!:��">�FY6�|����St�TV��"\w*P�(�Q�i-�{Jg�Ք8�S=��0]1��xb3�?&No�!TwP3�-�+���X�����iRxvƴ�u%]B��&�n-�Õ$c)c׻�fb�փƖ
nK�=�Z�0����d�tW:();45�������i/��,hl2 ��Ql7"z�f���jg&Ve�Fݼ�$��s�,V!�m3�I�!0?z !���&�bh9{��(&,�9z�����~��Λ����рyV;(
?�=�;m&��g����Af[vQ;���}ҽ�k4c�1}� �������T����a��v�M�qP���N��kj��������~*�9<���o^�8U����׹��`��?4�M,��ؙ^����>��L�"���]ĭv��.�=�[�m�g�-�mU�#�|hP��+��3��o?�8ft[$m*/�h4&��-�H�z6��)p�uS���|�V򋞖DG7a �)?�����Dw=��Iu�H{�M'��y�B>	Ի15[��[L��M��23  ��`?͊O���Ft�=�Us��k�����2�*���,
��ف��e/�)c�p�{�:Gܘ�3�B�	P��㑙:�V�ۯ:�p 6�ai��f��h�v$�ɠNXT;]���K$	��L+�����}@83K��L/�X��KՖ~����@�w?d_.(�C�D�G7i�����;��=O&��e5�-�����X�[�1.$��0꼒#�<[��8s��-��]���,�oWi�$�䨴aKmn,��.���$�li]���R%�Ԛ�������^2�� �M;�e�5���Q�-��ewS�^aKC�) ��= *���J�+9�>��	�J�6wG[[{�l��.�Z3�>6:�7^��Z9S�����mݻ��g�`�ՄN�.�L�Ŕ�ґjp�''βcZ#�8(�]�|k���DQ`���.)�������1g쀃���T֫�۪��o���=���l��}��L�T�\�8r
*���vz�Z��Z�*^ao��jz��0'U�EF�b"')��D%�!u��)�v}~͘���{�d
r��$���:ƗH!���F)� 9�N>�h���F�|O̯�$�|%���.������I�`г�h��N맿"u��8�!""$ �j��@��L�-��H��ɥ���S����v���� .=�G�X�]a3�z_��?	p��D �8��lSp�;�Λ�!�r|��V[��b�����/���:��A��ɍ����,������O��� ��uܖڰC��ͯBy
_g�n1a@U�m�bR�Z�d�f�Z*K�2�N�7�X��~�(�P��7h+�hQ8���^�O~r��ȶf�4�F�
Y걃���6��N
�8�$�t����ot_�^0#edȈ�D�5�7�dn;�)�i�6hZkhۭ�do�
M��l��Rش�u�w݇n��_�D���n��S@���vډ��3���ʨ%�a�1��_b`�po�n@@�&)ߺ���3��{YP��H"<ܪn��.�\t�h��?^A�\H-�J-��5��$߻�2�Ql�����ru���ɝ\��9zW)�$�#��#L�DEP�|��ﺑ��y�O��?a~$�"q>x]�}�J���V*�&����m|1�����S�<��rmr�S\c���'���IͲt6�w��s�D��鉺��$���Oַ�9�Qҡ��+�z"�d�����s4Ho2�~��&��<~1�E��bW"r�n?C$���Qk7�ݯ�����:��,W��)�&�d�"A��荧p2�f�bi�7���'�
ǖ�������&��\��-t�q��\���R�^���Ͱ��ئa���W��=����6���.ɒM���X}s���̾L���ݽ�\�HŢj�G^$��G�%T����g�i�dU®^0U�:�!��u�ʚ���N���f��+;��i��qq�k�?��>��c0ث�OlΩټ�#`)C�N��MpD( �����P�+ǻ*��e�
�mW����,`4�'ac^�f?I:dA��8�;���u;�l�b��V��H*���dW쭁�)�{Ot#�W�C�\�>�+�pb�n��K��,2]tk��c�u5���~|�b�S�U!����)36���p�I�������A�W#t��۵)&I`ڪ�.}�G�0=���	!a���2��Wc��R|��x�`��u�(��A�2I$U���vE|�R���M��o�.M�"&K���{�
�(c���AT-��q�����@"!�9��q#�Q(/<G������s�I�o�wǝ�`�EعZ��h�5���5Eo.�ڶ���s�`���&'��߉�Z�~l��Q��7	���.��znL���`Iɕ�]P����!���B~��,��	>�2E*��(�.�hy���:Ǆ-|~�)*44h+��)e�R\���DW'}߱c:+�ޓ5Gy�5fx�'�ơۨ�\v��1×拸ܰJĂ�����0T�EP�
 �k*�p�d���sw�u�_x�I2U�'&���N^*�B��3�P}!�j!^T��j�['ɮ�pJ�9`�.�g`����p��GH	h�[\�oA��1�A��T�7%�O��2s�uFd��2ƌDګ8Y�D�袀A�ا�n�E��Y�H��m��k����y'�&TMvh[Q�pl�͒��4��0�/�ѥc"�2k�� R���𥱺���h�/�|J��t����]0}VSP@:Z����~�y�C�;�exO[�w
K���<�)3T"<�ԋ���8䇔v��]��p�*WC�ZaJ�P��M�``3Y��T�TF�c� ��wM>�õTP��tL�:	=W��2.��K��W:��(.��_<�}2�Bn�P�����9`ׅ?�aOC..h��5C���I2�
��E7����H(�'�a^�f"�CՀ�!^#>�yϹ���R��7���I���^'l�����X�k,�yL"��iƛ���Rn�ڜFG����3�hr�/��7c���Kbf;���9a��qky�)�hK*2�um,	@p��^�l���M(eN.���k�_����?��QD�F�����8T��#^q'O���Z��8�U���E����"=�6P]/ί���R��H/����U��c���*��K|���l	��8����F���'-~��S�����v�oR+%�FĘS���aUK�34C��Ï=oO���U� e�_��
Bf*o|1Dk/.��vrx���|����Ώ���hi�ueȈVu"����1i(�p�`�ǵ��B����%Y4��4ھ�0a�f�"T �Oy�vW�Jġ�ט/B�Y��!B���;|01�ݿ-O4��tH���9}}BM�U�d�~�[��'�<Bۯ�b�F��I�n��o`'�K����2���[���t�8,�-~j����>���#�F��0ܴZ�߰C^2�kzL�"�r�^"I�nk��OF�h&�[��2��}Sح�#xD����hD�^2��<+��3H���KHz�5��?�Ҡ���ݍ������r�`ѓ2b�A�#�'��� ��5'I��O-���a#,t)e��Sx%�S��R���)�aD_t��
�P�<D��3��E�zr��G0���1'M<��d��g�����TN�7����4��S�ߖ�S+	�d�w�"�s���!e���v�I5�<�V,k��3{B"��K���?�.����>�ѸB��]=���c���>_�U$��!��UȒ�F1MG�̢{,ғM��j���@��I�5��Y�v
�[^��na��$4��GP�����K��FT�([���3�$����� x$���k�94��U�e�պ|I~u����<3\J[��$�f��s{r״Pu�^YO��K�;9@g=~3�$�Z���ϲ�*�W;!y�@�=��=�z��x��� )�Rg�N��n�M��֛���֋Rr��s;�M�X�M��'��<��'��G���W�9��}'�M�#���l�t?�� y���"^#V1(�g&�TU`O�O��� 3{�t!� Pq���Gd���/pU�N��,�d�$\r�������bT�wɹ�/�'ԋ�G�6)ڐ�!!^h�=��+�����^�飥�g��H�+�
��$	y�f�y�:`��gx��r�N2��T'�Z<Me�βS��1����]��~��}���،�9���v|�&���:��̢�����X�U�C�vr�@�0٫�6ߘaW��(��i�l���a'q}��D8(��)��5�/����tu�n.��5\Jc�|��I�Q�V�ڰ*�M�ܵ��!��/,;��͖|ë\b�KR��,	K�;��Ь���7�	k8^w!8诹9�����J5^ϴk�����	tM�w����Aѱ��I��t��e�aer&���跇�*�P�g����o@�Ƃm����{(NDv������(7�K��ׂLL#4�������3��w@��5������
��K2�����˅T�Q����*���Z d��
;Q�i��n��[�?}`�e����V��G`cv��|����|�˓�A�Xo��������n#	������l@i���4���V(���1� ��.Q4��&5:��eB�ڗ�S�F�ڠ�����`&���Q��梲�\L(j{�M�	���DǗ�|�uI�<f��I�@T������kd�*4SC��9
�G�e���F�[��U��c�$e�ȏ��6�w�R�U�U�|¥��D���=�/j8$����?QS0�z\8{.�������f�R:k�Y���p���XVi��hCn�Nq%b��<��M�ō>�֖�c䌑R�1���?�.���q�@��+��ܬ>��xRj9���ZV_�˸�#j��:�c-�Z��F����ck7o���� ��V�ub!���׹�����@^o&N6� �������]s�ߋ3��ڦ҂m���0��*;�w:��v�l��U���������8-hA�5ib�I(xJ����H:�ڛ���1)��=���<��!�����%{_�$N��e���ȖG�z�(3N0)Ujφ �j�t� ��t�A�H��4��X�V��FN��:V�&�#d�Q=����a���/�d�Ȥw�� -�).��'8�P�>�����'y�Og�u+|�b�-Nghm6km��(��F<M���i����<BL�(�q �I��u����XP{�XW���\d2�C:�Ofdkլn��G�%��	\ ��b%İu��i��sdڍ"�H��#淇�(�"�1���O������}�P�>Y�j�rn��^6`�W}�x�m�J!oyQ����2�fI�>��_�-|�#�z%V�a�"p9�{�x1X��}�@�2�Z5n�6�3O�����
"D�5P���)˧S�}�,{paJ��b���S�EP�u�BN@�����&�GE�8 �C�|�
 ok�����'M]����'N��l&wT/c��P��9�|���*���R7$;�y��j"�b5�5�{
tJK��n� ���P�1�>�N{!��C~��V�/��
TbOo��aʧic
o�@yK�`�Z��9/��� #�Jxw.�5J��f'}9���o��Ɍ�Ib`�6�S��}���bL��~	b����SBQ�~�S"��� ���s�e W&�h#p#�%b!P/փ�o�	��|V(�z����t"}y�����0W%�� A j�A\��Z�'Ȫ2���;F�>���#��Po��@�ޖ�<��RIp�d���)�]�p2�W!a���d�t&~���/����=�r�-9b$����#i`�ۏ"�3 T]<�v�����ew������J�����ȟ(���	��{o��(��F+,Չ����g���D�?���D*���-�v�l��b�6g�PK{�뚎�d�� �H`�)vA��Ji�Є�PUo���<x��Lmcpf�i�S�v^�ë-�Im����9�\���v%&	#,9� �H�UAeb�UP.�D�*ЀE������<�ҳ��	��N���锡���@(��d#�_�;�6�UP�Sy\L���V��U��������%=3�G ����'��������(�����_<Z�ft��?���Ѵ���8�����*Q����vG��h�L�m�Kޤ�F���;XH�E���y�]�P~�V����������Y�^�H�DN�[+QĪ�j#[��F̅�Q�{���X�3h�b���@Fսpn}�D�y#��l���m�LCf��eB1F�]��K͎�d	���������P��"��$��Τn���A6O�?{�9�b"��g���C�q1"�ޜ����(Ɠ�{���E�g��3$u����Fx��1:�	�FL�`'i���kk",8bHu�!���t�}�����^1�����������V_d��9
���ە��"�<ub
�z��䇳���v�಄L�
�"�e*I�ψ������HWn^���Y�(Cd�>"NW��l��|�>���ttʆ�C@�`QgZ��i�EU�us�h�H�k<�^ԔP���\�ߛk�Wv�{h��oWba�C��kYi�������F��;@ �/��|dW��/Q:�����<���{�!�
}e$�dΤ�F��M�� �A���
�B�6��~�T�*�≄��PkK��4�4mB/I l%#[����^��������Q��8�iN]����H>q=#H��ؓL���8	s	J��$ ��Q�-$r��lٞ�HL�O��.,��#�
�z��3�J��u�%{	�����qn/!�]��:T���}�+��H��t�\�섎��f[�<=��s^��Ub�]�|�O͏+�@<t��mk�7]�������	a�c]�D�+���%�M��=�Kڮ��X�5�����O�<P��jjsN�Z�`AZp�?;�p�	\&�:�ݮ�d�]~+�5��Z��sFB����Kҧ�'{��t]����˭ˑ���"N�����} ��:[��+<�R�[}Y�%qrAʀUk�K�U��ެ��5�pԓ��6� ��ފ�&H�a.��X���(#/t��@�\e8@I&�.�N�Z�2��ڦ�s˝�z���)��%�@c��PR�ctoߩ�Y���Ψ�p��AX����~�g|���;m]�ʧB@e���V��7m����qe=L	 ���hӁ�@��Z����ߙ�Z����&�jY(s�
��K8-�
�>��?|E�gK5m��H:��ۋGCn_?D�]�):��(��i0NٙT!���&�"���i�|T�3�S=ꜥK�1�M9{���Du�J~�$�^,2��
����>Bn�qB���1e�^�( 2wQ�5T�����D����T]<t���Qy�9=�;.�H�*V�9��KA���_��1�@�@G��3�w~�B�������F��J�7�;�I���N��y�w�L�[ȭ	sD���i�>�;���뿒��#@�*�0�,� � ,����#Ђ�z@��WZ�0�pg�5�������R�H�<���ec��;5�#н�iLn�t�&�4�/M'�qs�s�cVkC9'OGfE��k5>?qF����̋-�f���P���⿳N�W�;�tеK��.����+n�6,�ؤM�k�j�'o3��d��ʀ�+&M�4�+꿤��ާh���is=T���]�}V���]
X��4-A+ܱ����ʟ��b�z����i�����������D������t�@�˴H�AMk�k�w��Co��3a�c���꿾�p�(p
f�Y[0$3��҆N)�H<6>/���nz3��(|��r^������ux�&&��(�㸲۶Va�T^�1��ɐ��ip6����H�����ɍ���::GMs�EǦ��;�x�R�(Po�q��M�ϋDe	%�FB��+Q�;h)�C݉l���[i'5z�V�}Sf�2
���Jϑ�0-��`n�[#AM���L�Ќ�o���������W� �����>" 8b>��z��O

G��6�<}P`1�neg�����X�Ł�RU2[X�����J"��(N�`P�Κ�-�S��|kL*8���j���"��7c2�B��}Ҋ��$�#�5wn6�?��r���Z��CUo��Qo�޺���6�,nɜd%�i[)WL'�錹��?�f��"jȯ�:d4?��*� �1{=+K��{*�SCm(̉�t������{؛%���p :[γ2�%�W�̽�)����$aȳ)SdD���q�&� �<����t���ŕ�e���ΛUA ���aa��hS]x�>iJ�����c�{'��]T-���AпnIWT�}��D����2]���@�uq2pp��˄���cҔ9k������6ij��-�28Q�n�Z�#��
:���Gx���W�5�����p��c��Dn%���S#�H���BH����.R��rS��{1�{g�j���\V[�:z�Y������)H���/|���]���)]V���/)����EVv�IJ)U�~K5 (Us;���!/1��B�O�z��=�=�X���,g��dG<�o�h��q��� �,��)%s�P4�,���7	�f�'�.a��Hi̭8��'�f�\M.�N�LI�5Ӗ���Ù���F(UU6��Ii�m�h��Z�A2.U@�9���j�!9�i�CB��wJ^=:ӱ*��T���P��#�����:+���0�����l���(f���m[AѮ21��Y�1�������P�W�����tm�G��r֔�K$���u=m�O&���&o�CW����W-�����$-�uL�`UM���@�l���b����0>�ů�UF��DⴘO
�E��hst���q�e��o���Dt]�I��a�D *��)0F\c����c����{�A�V���� �?Zg��ƥ���ERwcr׳���}�� �"��R��ΰ<���qy����[߫<9���5�`�����p��S|�\l�LE�q �Y���uNg
*h�|׷?d������
!�w7�G����f2���X�v����M��%J�c���u�.��?|]��k��*��T�67υl�(��:�p1�]��>f���#�\�EႦ�p[� ���OS�����R�_6����7܂?�3��ܕ�PQ��n�"AĕY��E�c����c�h��I�d�e:ɋz��{��m(��g��JwX�E�S�d1=�Ъn��bLr����'��D��.���8ҲJ����:�{�{-�C�=�_љ��N�80�`?gtF�_�u� �U�9µ����Y6��%�~MVW/?gw|+�BQ�C���8�-�ͱ��&�{(�����J�����RE�G�Z�r}��<-�X�5��|ǍS�v�S��O��᷺@�e3`Xq��t���6��o7#¾�x�9y�6ѯ��%����g�j8��}�Y���F�(�q��l'
���ry)��1�<f���E�.��*$�Y��߰�8&� �R.pO��2%�����֖)?\8P�r�%�I;��eGYTs����fX���Bܱ�y{�h��'o�_�P�N6P<��{#d"/5v�&�ڌ�؋?��Cs���je��i#�E�k�[�h��]���:.R.S��_�G���3 K+>�$�Pn�-5��cϢ�^t���=�}�׫\��<!)�g7{����b�ޒ���9�?A:�o�����Y�t	y'�)+�`�aƠ)� �9,��VdeҼ��;���TT�[��������-���c?�,����V}#>O_hN.�=�K5���g=��o�緝�z�r?;,W,Q)�B�E#o�EgM=��S��i�Մ`�z�����+��p��|.j�����0��Vǆ�::�ͼA�$2�՟D#a�d���'�~P<���D�
~Ǎ�֜��H���H�T� ��CZ��Ă��6��C���'~�CSN)su���-��������V��30�V�X`���v����l��3r5�8'8�y��sq\���$�W˥�Xmz��MN��Ҙ������+�%>u�g,|�	1v����	���F�l��A3v�Ӌ�K4�*��jJv����=c!�DZM0:l�E,�e�0`�v�X�:�J�a��y՗g���'4M˭�F-�v�dxu���v�3�=6��u/�<��)�pD�}`��}#���a{��s\����x(-�.;�GsA3j�y���S5 2v�$6��un�=�qDXx`� �W=���ks�A�����}%3o�f�ݰ�gǍ;y���8�f�H�Z�+�G<{>�4[L�kw�:tr��,�:�{� ���BfX8��@Euŕ��Vמ
\�o���i��_I�JfS���b����?�q}G�p��i�9�_�!:��A_P �w�#B>T(ѷ$��Vى猈�%���t�|a*.�8�f�<������#��Lk��Y�j~`��!d�y�;��m4�Z��"R�u ��!V�H���sŕ���p���݂A�K�
�>9���6ר��1.���c��͔�5�G.�n�S��m��Zv����:�U�T"{�K*̹M�g�����f#N�,&5J��E����h˺Ŵ�:���줒 �e��.p�$SK�k�M�&+i6b���/!!.l[uZ(��@��A�wG����ئy�Q �V�cm��[�X2n� 0�wdw�ijv	�d��/m���"4#�M��L�џ��21y��MY���j�
Z�]����6AY�H��^R�D�����Ҝ�f(�#D�����7���I���v���!��>mD�5����,8D�����LZ3	pI9�O�+|�
}�)B�3{�����V������=�4h��[[�j���{��׶J+>����ѳ\?�U��h�Wx�T/m|S��BWxA�B_�T������5e�eJ�z������ubzM{����Q��i�.E+�xP�4���7c*�Gp������ee{e���QO��:�F&�B�r>�Opq����E:B�9�O��!?.�2�A��m�6&O�� t�_�+Z��s�����3�9����/��K�2�dXqM��J��]�\���o�L��p�tF9^X�G�;J �YlJ�g�cǸ/�C��:��(��fz���mX�n摲n�I/�)_�������8鍛U��@�`���&��z��Z�\"1�Х}b*���T_Z��2^�y�Zx���Ų|U��~�� ���`���TlX��(\Ϳ���AV�ĝ�`ɀ�o#��H�t�~�}����b�3/�f�R:� �ϓc��"O����	��D��8��ͯ��	�^L<Qo�X�~F@�P�	�S$i2d�l���:�u�^�(��$�*��#�9ھr�B��)���{>*b��y?�P��6���z�y7TI��[������K-��Lvsm~�M20�B++a�`��������f�3�xϼ<{�p�7���R��2�K8~"����"t��Z��
�O����(3,Z��W3/ ��󓤖Q�!�ؚ���	�����mr$T����=]p�'pY�&��E�[���=<:zD���c�4�"Hw˕v�5[�4�Q}J�]_h�d<�r h�~���)	k�i����a��~B:�ENƐID��h^��N�Z(����Zg�� ���j���6�L͑������A���n� Bu�N�o�s�D*�س���S6~ ^Z�]R�B�=����ot!����(��2hG�R 	:�'�t�!�$�eB�g(D�dԤ��51�խ�0�����h7�NI*:_���6ڲ 9Y��J2-��+�Z�I�����5�E�����o�Jҩ���^�K%�'T]���	��d*.t�.B�7_��>XE��I.Y�Z��#�Y$bggJ�RwhB�ό��)s5���mlE�W��Q7Cr-�TK��ﴨ�N$�^_�y�ЅZ_�o�@�J[:�aP�l��o@H�l0����}@�Nù�C^C�����KO|݈�#������M�\Ԭ]�m���{� q?����PЫӶ�˥�K���O���Re���)	���"�G'���Iy�@��dWc�s�pP�h���#
n���,ˍ�|�P�	b2��t�0�F�eVLO'�����ę�o����]�w�
������ѿwe:%��۴�Al�`r�e��`T�M���-�)���y8���(���U�/��1}+ה��"�~�pN��x�Fꗮ5���a~���'�����8�G'��me��.�ʆМ��3�N��ҙ���W�ӻ�`�e�f����[��ڵYᄎC�P��`x2q�,����U7K��WHɿ�ao�Ж�X�:/�]	����N��Ƒ���A�6�<Y���=#�6��}���[��k��C��!�}������(�@�$�ܴ�����׷ �}��hdѰ�I2����=���aU+A����،�V��÷��|������z��I}
(^a���uiVp�xY3,��7h��4���?�yF�J3���1�K�˥ ���%_	5�(�{<��o��F���e[���*�h1R%�4��������~��i����!TR��>J��4�:M,���-;�H��&�z=�(ǚ���D��ʱِ@�$|�X�������{j�s���d�2�G����X�C,TԛL��=H��;��C��;����5-p�S~B�|�����TT�]�<�C������GW]��|��������o�8���e=X��r��Vq�j���N��}��}��[M�=Z��g��e���^]s/���c��0��%�a�L|��"c�p��k�Qbn*`���_�	m�b"�^3��(',D	�ȱ�a���u��2e�ݐ��@}���2�F]��w�X���EK7�v/'*��v��ɥn7��1-촷�xr*-t�2�VA+֐/��b��L�;��^,�V��?�;��f�/$j�^C��*��峱���LK���0c;���Y:�=�}�/��v���<[���"�B�<yLD���i.���*�+�f�J�-bHOm�\��~���f����򌗒6<�e�-�	���P���آf�O���^cUl�N���H�i������m�-P�ţzݸ[������ш���J�U�2G{�K�'.�����j֥���u��ʗ�q�\F?��H�����|L��7�X3���_«�,�_`LmM����@������&Iv�)XQ<To�dڳ �b��0"N� ���ѧp�w7K�I�P�ʻ��|ifޓ
�Oh�ƻGJ��5r�r���1<jP1��/��8�0k��/�Ƥ���t��t@f3�5Q�xv�R�� ��H��߆WklPM�m��0��~'QF����7Ԝ*���K5�w��s��Pr-Z04�^%ʄI��Р�<��*ae�&��g��<%��䉹��u:;:d<!R��(�6����7�	�C����J��hZ֐�_I��6)�dC�~<�&n"������EG[Tihj'@?�zG'�2a����?�kA�����n}�pOӡV: `���ܾ��-J5T J���3�����tRI��k���0�/�����d*��%!P�g�
�R|��g��S�)�0R���ς�5��@�Y��Pfl�������Y;�KP�#��$W'�-SU�5G���JC�}�+'���`c�@pLV�<L#�$R�������f�D�\?�C0V�˸����ӂ�W(WփMkw�0g�9f��)��i$�Ffu, p�д}�0a�4-3����WBn�����ޯA���N��mI���߆ßԳ4cѼǯ���C=��\R���h���T�s4�0�D��C'GA�o��z	!�����=}����;�C�zP_1l< �ipY�*:h�����Baw�Ǧt�<}7�$GɠuĪ+a*�{��#&ݧ3�M�()�4KM~4@p��g�Q������欥��A�5���:�Y&����n��[HҔc����͞ˡ@���19[vQ[���������ݬ�{�&�0�q��4�
r���V�z ��qQ NL�(�#z)J���C��l�p��q�e�*��aU\S��ݖW��1[A�z��QAD�a�[{j��l��(2�b$\h��`�o�@Pf���8[�C�G@�܋{lW[��4�q뇆BMIgΓbl^ݽ���u�ꌲ�p��R%3S�I�^E�{�*�4�MR/+S2Y4]�rl�r��Ĩ��:�yz��pEvt�rG�U��ւ�I������R���%^^�@m��uP/��A�F�h5P�����:��Jw����P����9�b���i�E���4Q���QN�(c��i
�4ud`���u��ĞL:m��>X�L7s{5Y�I2x��+�xȍ9O7i���
�J!v;��=�<t�Ϸæ�Uɛ�w�1�\�z�J��g�B�@�֒���tB]�0�$f��O�mC��0e�F���>�7b��f�9L��x��K�'���{�p9T��X}�@�����D5�/��G�tZ4%��[��5O�g��/�滴��.�@%�.�Y���� ����s��,f��J��v�!?DG�)�����WB`�Z9�ӥ<-��[8s"����#�����K$T!��1%��)�V=e��j�W>���>4	�Ͻ��/S��]0ag;c��6�֒�X��o��U���"F�((~���0��ş��iP����Q��W�Y�n3�!k�Zy�{�2#
S{hͫ��c������F��,�I�N��]c�]�Mؘ9R/W�)W��9��fA�0,�L% 
�V�魎(�t�{�J
2$�q_�������>O�0�n���g��/�fw�t����x�u���3��hh�Mg���N�i�Y�"����+#��inU6;mF���X��`�m���W�g3��dO/�'t�g�Sy��M���,|c�ّ�ܰ�5)BQޖ(/���l�����,S?ۋǓEХ���kiE�~���fF1��������h��ެa��Ⱥ��X&P�9�Ι�k�յ���1/�)K��h]��g���P(Q�0�o_�q]P�����&~�do���g�?�ƤPT�&�({��fS6��l�?{���V���B��-m����p�w<�Xc%g�e�#RN��3o�w vGs~;Cߗ�5�6c��2�B��"콨K@RE�ǒb7�sY�-t"�.�T����(�u��8rJw����A,M�ɝ�09��ϑ̎.7���[h�k�mPJ��É�3&{^谷�!�{������;���B��A��D�%�����/E�A�/Π�h���.E'"�Xךt��YK8�zG4�@$h����!خ��-��E���K=�_�:g4��qo1�������fOdRP��h
T��>o@2�Nb���t%qf<Jt��D=M�"5n[^���x��Y������G),�^�D�~�.|W��$2�^���K��d�S�)��:�a�&&�έ��mIdV�� JJTe��h�6о*���a L�b�?̤�ij��ۢ���ߵ��p�KJ7["���/G�lr�/��@]��&R�J�f����0`��2�sz�=-RTȿ�.a�;��e���\�({,�sq{�����z��g��5�^-G��}O���9Vrr�Ͱ|�Fq`���.�P>y���Oh��i��
N��ޯ�Zh ��^��6�?�Bǋ�؉0�;ԟ5r�,��;�T�"D?"�`r�Q�ۡ�08�K��`MQ����V|UN7��(/�V�D�?r���Ub�+���'�[����u+�S}��Ӧ{M�5�m�J�
��i���a/� ���;��Tg9��/���4}�9ї�=\�"W�]��aGq#�d�9Z{�
��ILf|e
&�;� !������ �u��?��&1���_�<���V�.���"�W��ݱ���/K�,(M+��=?�<��_�җ��������e�=�#��7R�;�x<�/�<���2�hTd:w��Ӑ��ߕf�m;"|��O��x�ʉ� �O�<������Dt_u�Q_J�[BH/�z�S��#_=��wڂJo�N��DpUۨ�����&���o����A��'�J��S�H�9�E=�H��k��#\��t��+G>�}�^+���v�G��X��c�K�Lt<=�@ ��8'7�	J�]Ĭ���M��=�ϓ|疿��/��ˤ��Q{�ܓW�܀�
?�\�[E�:�C�w���0u=�:	V$Y hƅUx���^RƩF����G�@Z��T�,����Avcm�ph"���z��5 2K�A�
��D�3ο���ʝ4޾b�8����֏�q���Ӧ�e����]� Z�X{b�m�q���fm/�� \Z|���}��TZyt>�}�}�݃:]�����Y�Y�2;��U�0�4e�A�����)du6���Z�KU����f��oӕD̆�$2)�3�:az݉V�ʋĲ+�V������'=��Qis����H��PҧZ
şK[	�-�ۉ���%ͩ'_��xh�WaӉ���rKS��h������}��N �I�_�&Y�l�,jl.x#���7��& ~�8�|�rwG��(�+�֨z�R�{��c�κe�]|��q�w׵Q�q�׫Io{D1e�C�JƶdTA�(���R%���8�%?�u�uC9<M��fL6�PP5B����K]����#r32]����T�fs|s��7u5�@C��Bw\��ԛ_����ZN3D�����O>T��*�{�9ʩ�8�1AK�8�f�� ���aG�U\��+�0�s�����@�\�}���9����L"p�Wc|R�h ��s2
[�fz���Ԗ�'לC�z�
Ro��#��u����4��Z8ְL/-m�f(+�4��J�6껔��U�m-6����Q�tѪs�xO:,~�� a���)!��W	��;�
�Ԓ�FY��¶��'s������ޫE����|�`	��S��k�Ͼy���g�?FT	����9#p�m�G*	̳����Fn��A��f�XcZ���t���a���w.fa1�!���"����:� ~���ͿN�S��9����Y1m���dk���;D<(���U���P����6r�%f=�AuE+�ݝ�Y��������/$�J}P&�y�`n����k�Ľ��r˛^Ғ+��ؖh�p��5�P)W ~����� rh�b���Y�m��8�hc�ߚ�>r�5�����ߵ �4��d�F����#�UӢ�Yn.?e�%��!x#l��)�>��j��K�eQ����A[�r�G\��8��$J�Ǚ@����E�˞\��p��<������]9�c)v�Qx��̊�p��^x��!e�D7@�"9�� �K(�����0�M ��7ݰ�K�}�-�xj5s����@w��!�u��3�����܏��kU�q�Z9�Z[O5�+��%�3����������q
$|I>$���f`��]���!4�T��"T�ѧ����Zה����RR/�#��OB���IRFC��Q����oZ��fM0�# y[qz�dE���biS�Q1�f\���_���꩓k�G�'���
���N��Ի!'ɧ�ЖBW$��C;�`�.�����qJ-ѽ��|�g�uCZ8d�`D������;=�X�;9[� q�k]o��I��b֮m㣃	���ԱĆ��ܗ�ȟ��?D<��^��{�y ��C�ti+#T�Ä�_-�=��2;��x8n뻠ĩ�{�I�ë�=����=�VM�y؜ÆP���3�r>j���*,���Ē}=��P��`��p&�j������k̵Zg̦�6���9�%��G�>f�/��m�`� �a�F�c�҄Ž�u��K�[�X��ɣ�	�����*i��_����1�n�5GtBMP�c����H��[U��e5I���}@4������\Iy���C%�zR �hDq�>��;�����pn���Ybxos��xr9?x�����#�-�� ���2d�l
�K��s�I�|���R�-2���Vk��reJ�DB<Qt(�۠`I�XXNN��UE&�b��{�6�1?0%VH��׮�NS3u��N`,�l�x��s��7��q/��Ur���	xU,PLj^�Nk�[R�L���~n�9�#ݖÈ8�&V��U5��´7+T�mQ$���n�;�g���ť|��]�v�J�¼$|e瓼��?�̛�l�+넎rK����Y���)'����0`0MnV������� #�p��G<�f&�9�"/]kEc ���{�à7r,�K^�׋�!�}~��S��9⺦]��5''�n���r���t�|@��,��M��n�I�
����6n�2S�����qrkB���Fc|u(��A�rw�����栆���3�ۣ* �z��1�H�����<S&�:B����v&3Il�Uxrs����`�~K2��SL7��WGƝ%�ǔ�KX	ǭ"ˠSQ.$�V��B���f2\�B�9�kg�O~��`L%?�MH��5��OxVt:6���u`���4(����e���jB�f���R���'Kť�݆����z1ջ�k���(x@��/4�t�ZYK�Ԣ���I�A-IT��J�FJ�pr!���`U���"��Ȣ��Н�_�����0�2\Kc���b��Q�$�uS05E7Ǭ�	�`:���\K�Y���I�Ɔ�k^�� 1{�W{;��
>eg�,�d6�dљN�?I����2ײ�yZ���@A%+�W0���+�zr#f�Fc/�0�m��˦{Ώ�+��2��o5�ߣ
\��:i�����ɓ�UD�)ǌ������B�6E0������0��!m�W]l^�B ����˼\�'�^��7g�+�n��D�y)�2]CP�,��v�벋B��!��JG���,�t2�����\���]�����A��U�A;:���؞&ok~Q! ��L���n��������!K?� ��j���6���.وXsq>���ڜ.�S�z!�E4�#��<�Tƹ�
��NL�O�2����b|'<��͠���,���f����u��_��l>��Fb �N�Mp����*0A]�q�u�q�å0�9�%*%�1��G�C�*�j6)�")4,va驷�iDӵ�}MT?�T�z)���8V`Յ��{Qp�pn��KhNȺ�H�V��A����t��ME-³*��"1����ц][�Ò<T�n7�f��R�3X,��I�D7�0�0�.	��B �0������e1=;�]M����#��a~5�6۾rJ�R��ә�����5BY�D��McO�����%,����Q���^}�v�Z
U���
Z%���ЅI%~X�.����Y�^��~�!6b7Ԡ`�=�6�g"k�>�Du�4��f*�+r*{�O&�s�mn��Y6-n��UB���pFζK�u~b�C�7�z��n.؜��t�>ri������t��Ṡ9��b��������'e�X�.ޜ��SX���	f�n��j��aT#�Ǥ�ǲ��`���e�ptȿ��CL�ѬŢ���-�-Ț�q0��'#��Jq�%R�$��q$+̲Jdh�r�a���b"J�'��`�i��#�D!q�8���:�=!�TMj[#]ç�u��9~�KQ��N�d��eA�w�M:G�Q4��-6�����l%M6�,���"�B�����t�Z>G�^��@�Jp�wk�H��S�*���Q��5�o�0����'�Ɖ�C3�ǞD�Id�V��4ŊlM������:��=�o<�ȕ�<�k_t|�>q��t�0¦:���\�o|�:^dW��mV`j���@�r�pa���D�W��h�H��c�HJ��Ֆ��y(�!U���zd֯?N�)����'�MUӶ������k��~�E�u�z0�M��3z�{�}��C��m����
*s͟��:���u-;D�p�D*�S94��j�Yv��;�p�L'x�^�6���[� 郰r_���c
Qa�'XX�L+�D7g/�B�����3r����SH��N?@���H�(��N5��X1����|	K-r�=`j~���_�O}�0��i����i<����1������n8[�+��+�f7�GbO����5K@���7������yF��"C�b/-wę�3�r�SAs�
k��k���g��ޝ>��,��}�
< ��5��k���}M&l��U.r���|�&�Z7`���w�����T�W����+2\�Y�Y������3�����d'`�(.U�i���h�g>_���*�)�B���!:(�AZQ`
�4N�M���˄�����<���à{p�k�q��K��N�dv�>Ș��r�5�zX��!���J#���ݐ�
ä>���(L	�h):7\z�M��oU;�����?�F����`�ОQ��m#�}��Y�3�0��0�����DR��
�g��_��Aè����%/9�n_鮪|FOQP��:���xNLP	Zt���d*�3�œ��l����7���Tm�/���n�a�����_�����h�YG\6�ǧ<�S�w��&4�VW��ըȼ����xm��a���d|��P��h���Mu��LT[3�G��y�X�ߧ=؝�(���lKYI*�����?�����u�M�\�D� S �mՓgf�v�Z�Q����i4
_��Ds�Ωx���=3z�����qu�"�S:���ܚ���w�����l����K%�Z�-Hގ���VG�h���}��y���o*L�\tRN��[�1����o�^j�.�M�5���(zd��%�'��`���Ұ6)�"x�5ezC�\i�R����'��?���~�2ꊴ���N�1T�R�D��)�n�h��dT�glͩO��l��>�� X%����tV'��k��E��6eg+����쨓)s1�EQ��KG��l��~㽧�*�ߑ��b���5.�2�8IQ��9K�=2�S����LC�o�PS*�����A�ۈ���N�׀ 0�7�����M��]�L��+�����w���(�9O�Щ�	Lׁ��zW� ����j)�Q'TUpی�]�Hty	�ZJJ�/*~բ�9����h�k�	J�1h�:$��`��%A'��_O�ç����]+��3{_y7)�)�����ro�`��ot~*S��KP��\��aT6-C"c�����¿� ��T��"M�+H�Z�x���%0��@g���92b������{?�\���8��F�D�
 ���i*��]�+�C��V�!n!��j��Q�Anj�m[h�eH�=�< ��K��^+�����p~.i,!6�!��e��{.���&�5|	1���1�(2����HL�[���Cǧ8:�~p�Fk�`�8s��]�E#߻���t.�Vժ:a���/��] J�E�Na�m�ֲ�#���"��n���A�.���p��Dk��s;���C��L7w�d{Dd���B���/��:_����\pۏ�b�,_�����!I*�C���{���.�������_$�����^/���K|/ى�	 �k�aD�	7%!�H���Bu��rZ��k[#͵J9�(Y�����k4ԃeb[�����n<��(zI���T����祶*f �t��ԩN=�|��%��Y%_����S3my	|`4D�X_�<��8�I�j�����gL��OgD��ݾ�F��4�ƛ�uk�M-@d���H�eW܃U|�i���)�Yf�	��0��n�S����Y�*u?!DY���9�T�Ǌ O۷S�^}�<�ÿ1���vg~���w�4�UЩ�iA�m�U��*A�g����_�Y=-��1ʬN�F=��R����~�է;�	l�0<��͈�2����_��f	X�e��c!��L�j=7:����x^A>����7+E�#�~/<o�R0�QV�+��]���ܨ ���y߽J�^x���������s���h0�[��$J���Y�w��zxI��./��^)w����[�?y���3��QP��nB;�K	wj+1�0��+����^�̟�䲆y�.w��00Ǽ��PL��6�{G�a �SG�Y����\��yt�r��ϯ[�-,��X8�������S\g�_����'C���k�۹5��j:�M�����}(�&�m-�ѡ˚ �0\`p����`NL%����Yѝ��qn�d���3�6�׀.��hBE���i?�G�u2��>璿� b�T�8�>����<t�5��|��H��r2�d�+�H}� ���5�'2��U�E3�'��X3���m�}�z��>21k<]b,bȻ낻�x^ψ��=uh�7��b��Z�ف��M�B�^����O����A�q)n%%��X��.�1���}�������-j<���I�� ���%S����Û~��e���NΕ��01;�Iv#�pڹ-��J����5���-(^BW�>{09����O��g�{�|�+�!���;6����(|o��: ���G$�K��*o�Z��w`'���,b<-�(�Į����Z6���8_��%؞�)(B�6(޵��Ӓ��r����{F�:(Sk�ȺVLX8ad:��0L!�o� ��Xt��1��A뗊+iwcU�g��M=9��0WLT�A�<6P����i] sz����s��hk`6CJ��Q<�m\�8H wn�̾P��S���xgŻԢ[�����S�#��uM��W֝���ZO����ַ�9m��C��4�4	1�L��w�zN�7�ݩ@�����s��L���:��N�>���Y�F�a'p�*��7�@|�x��9{xٯ��TO�z��l��{���S]�*3�x�����[ϗo547IO͗��^��/����F��>'��Y�ޣ[��5�M��i��;m�6"��:co�ͫ�욫���y�ӫ_��։��P�.�����O��L����'��rT�d�#c��M�wy4!w-�N��f��y����P�t�����;����/=�h
�qq���)x�I)�N'v�##� ;p|��7&)m�č�҇�M��V(����R�p��z�L#����C�8Om�r�r�O�n�?_����?Ӑ���MI�z@	�2��):}p\���l�x}�	�w�H�贝u
<ԭ0Eg��=Z�R����tw��Z��w��F�=3��^�#~����-����:��I,�J�0��Ee/g�B�l�m�c��q�ڳp���iξ��S��xPEϗ����u0�J�����(���5�oف�ۥ�-���N�Bc��4�Q<"sJ%���W�-T�gx�M�%G	�!5G4�Rƹ.�D�O�;�d��	���Gp�M�Ԑs8��oՊ7��v�:Dݱ��{�Av$�$Y�]�&e�L�A�h�W�)����R�m�}⼰ T3�T�� `)��neTc^�c�愌�Q�����C��P=�s͕?�U�<���'|�Z�����54쮗ۚ� |Y�����O�̩!�Q�+i�<>�E�[�����g=if�|#��%fP�~�ޞh-�>"���:e�AFRc�c�v>�y6�ʞ��δ�3���f�Z�k�(FPN��|_���z�Q3>�`ᓶl��H��A(Xb�Kl?i(��M���K���oQ��*z	�,��_ĢUG�ְė�;5�[�7�2d6Ո��	�
��CPަp�HX�=m���5���)��>E7#�r�h��:{�Yo�ʓC�Ţ����<�Ug�V���H�p�y�����d~��#��jq�MA|�	��,���tj���t��	Y��	�;\)�+�"7��^�PH��I��J�B��}�ȠOOF�x�ǳ���'a��=ﺲ���� ��y�Đ-3�y�&�k�5��^��!�N��/���5��<�7�F� �_qm6ԯ����zG��\4�B��3e$���P�H����-PY
w�D]��A�1���J���Ȼ?Ƽ��භ�l=�M�IS�X�Y���Ldb~�i�a9�.��F��Mp�����v��8G�~p,v���K��Uq��\�ƃ��}����A�I�M�K�ɫ���&�9@R�}����п��{1��Y��\Xn8�l���E7j��:�v�
�����PsCB4�=�,�&����/=m���K��"�NPG|o����9�|�
ZO����o�T=k�)H��m�d B9�ݱ���;<�G�}��+�$9�m��I��7�P2��eݟ�E �U��VdA�&�z��7��O��}�S���1Q% � �e��;:�C��n��m��s��l[�Eߕ� |A)c5.��������&kc� �b�L�e��B��%���,>��SIJS%��|���3�f�vcDˮI$�`[�c=���s%�Hp�f�s��6W���-t
_/x���hv-���^�� lktui2�P�1���F�1�'#��kH�jo&����Ei,z�dV�^����g<�l .�mB2�잨�E�"�I���lWD*4���y�����39v�u��G��G���"�_�������m�W�u��	C�Y������R�ى-��0���ȷdh��(@D���Ԙ����x����ރ��Ρ��#��*��yTK�������(N\]z�"��7��]�oM�`P���k�����
x,Be6�V�ńN�?�mMr��[�����3|Dbb�j�]�|'R��/T[��9�'2g��Pu
$����b��bv�#Y��	�b�7Y�]
�������U`���>�k���CK���u\"�|����P�4]�[/`\Y���'�SԼ+D�N^���XNL���%$�a�|qż���ÃP�OW�_ʚ�����vTL��|B��qi7�6��.����
?�k�;6 D���6�C ���`%�g��Y���^�rx/����WS�
�M-b��pKF.Pj��,�Ʃ$����O��ݽ���*Hv�)��z��v����5W)���_h���s����Lƍ+����H�P`u.��k�0D�@Ҏ8���%:$�Ö�� ��t��Wz�mgK��kz��$���Ǿ��>��c�qD��w�<�@H�jO�W�Q�ηO�U��8�-ݓ�̌�C�����xN�)���N������e�w�GT��K~O��ɒv�b�}7Tu����5+��_Q]�/�@ q���������H��aN�چ_Qb��Q��T����"�0[Ze����Mܐ�wx��#"������6��LHM�� 7��լ���
�Z�%��r���Ev��E���CD_L+�8mqH�^�e��DgP��R^�.\W�z5�;� �w!� �����#E�
��W�nı��&���j2���/�hjp{z]E�ꏙq֡c
i"����c����r*W��{�x�]���'���^�l�EqG����wُ�H�<�� #�E�~G'�Oj���g*�˭�%w°�	 Ì�5��6B8g��&��������t>o�����Z�w)���'����d�%� ,��~��oh�y
:�M�Wh�W�����{EP����n@B!�p�/���Ȩn���C{"�%8�5��;_
���޵K[Pv��X���՝�ËX̼�I�W�f}Uvt��@\fκ_���&��^�~L�$�7��JѝB��P���Y[��Fɏ�9Ij�{"�yԭ��3%�q�=�S�t!F�_��@�X�)Toծ�/�em���J�of�5��i�i�1����nR�;�t�� �E�{g7��T�1�nU"��^���!W�\QT�39�n#�����������+�M�4r�K&�>�	��"虀ՊU^�g�C�Y��Z	���W#�o`'A��_�d�cF�{�WL�X�v���,��m�MyjĦ�k� sl�(�*e��x�sý!0��P���ô�p+l�	G�=o%���o���&�)�)Z\A�N�g�߷�=gO^�Eř�lJ���LQs,��>.oŒ���w�Oh
���/�י�{�u�u\�t�@hܤN)��vM�Q��)�'ө��5$����D�8%lsO"���*">���x����bC��p����B�:��R:�J��i٧4h��4������ɧ�PyW���()�TQ���F�3��V�]r)0O��RQ-�!^�V�9§5�o����F4?͉c�^�&���J/�W[5 Ts���;��ds��l�鷊I90��4�kP�.�S�hâM�x}�r�L�&l��>����<[�����+�-/�_�C�\����ӣ�hg� i�4�5^=��c]&�ݻv�F� wd��skc��O��%8O�5%P`���
n�S۟ɡz�[șneP~�R�,mg�jҘ����z�N��E��Q��Y�!����	`�I��}�tc�]�պSX��W~�[�k/Df}�y#�3L��W;�5i����d*������ɯZl��r@�p .��5N��(��AN�޴M��WaJ��b����VɁԭ=1���-���Y���PIV�z���j(�#�\��Z��!��_I"^FTE�������oի�=��С��ōS�۰���4 k��-���f��Z�SʃǗ����
�4H����
̧��)���i;���>}S�~\�U�<:,�w�F[o�z	���Q�
��.!�%Gg��-�� ?���Bk�?2�)�9�4a� �}�>$��p����Q��F)�8'�s��:�_q|��f�P���`�L�!9	���s���V�$����i�[��S��ɰU�~�.5��Ό6h��][^3G�8=�7����*�ji%��O?�'���o�t�׺e�_^ͩGa7�}�o���1��ƭ~�
(�v�HR�)�o��y�=�ɡ^`�UT#F���l���F(��]8
@� 4�}u ��q#�l���]^b<KĊ�t��WK8��ռ�)>���)�9�(^P��G�X��ﱼE<B{@%�ׅ��8��<b�yTՕ����[���7��C�M2�"��gE��$��LG��~�cDZ.\7I��U Y�΂�#��K핒�L2��y��1�#r���X��=��pD��Apm4ꢊ/��o;�wfH��|�N��s�)�h��4QZ�۳8C��"�Q�dH8�ƾ�[d#D����`��yz٘S�A{d�qH~�7 �D���}v�j�&�����]�E�$_&�&�:9�6^^����������nͮ�}xޗm�
�7�C�=
@M�"w �ڠw���1�;��k9�R4����{]�+�UR	-l��P��.(�sba��x���k����1�t���Q�<��=���0s��GА-*��7b�}f�j��c9S�Y{�"af�}�[LK)�C��i�{k�~q��j&I��r
{ˬ�/Ue�{tq/�.S�fwI7wl�{R�3l��������Bǆ<?w��A��
/&@��(2��+$����^mR� ����f�*���Ţ����A�$���<1��(�)��)�J����9���FN�-��Tr>�2.���{��!���8�	�U�f+Z0\}n�7]��[��`�C��M$�>a��pH�u�L�6QY��Nj`G����w_��!��=/����1�zZZ��a�s�GG_�!0���L��o�hiH�0뼈��"B$�K�Y$Ztn�-	8�L����w"�C:���u0e��ٮG�ؚ5f���P�Vأ�1@Qy�5� Qv1�P�����$�≎��+W���iD�S�r�#�s_k�n�.�X[;{�\��&W�:E��R���f���V0!vX�'p�����l�Vo�7�$:>����H+�^��F-��%1�ܿ�(	�_���괍G6��c���U�^� �����b�u?
ٸ��mh%kpC�q�?��i���	8I��1��Ҫ��U�7�1����񚀶h��Uݐ4�V>���'���W9��F�#���Ջ�H͉8&�˯A�*̎�lk.7{�����0�������՞t��<�j=[����vHҗe %1����� wt�:��%�^�˶����B~���	�)�s��#{AHׯi��,��$O�#������u�|�Ah�7�q�:��&�0>f~^C�yK$.����=�K�u�N��k�{H���n���1��?S��Q�>z��Up_��/�< �F��e"ov1�����Ge��nE&��@��ׇ��x#�BS���b�v�l����v#��H�Q5��L�����N����Xai2�l���	��j�ud.ǛH,�eܣt]<���"W�=�U�@����3�6Ä�n��� %H��/�:�^�8g;�E�@j���h�4��H5n���}�R��b�Df����,��]*vQ�kZٕ�&�SE�m��!!��R��1dFX3�ID�,-�.ANZ�$�Sԛ� �j��T��=�Rg��MǙ<G:��\C�$~̋�t�DŬt���!h�O%{(t��%f���ѓqY�Ba��4\Д�Ҥ"u	@]rB����tx>�:6�����>��*0����Y����R,RnD:�$Cs���૚�
��(wPyo�q�{\�6�(��0+}�EgAe��K(�#�1f�ji<�&U ���+IQ��s�+��8�2�K��V*�\����A�@��mnI�q���s�A����@���-���ۥ�7:t�cأe�*�o�B��s��΍��ߦ��ç�+��Y׻n馫t��-��f���G���]��|��͋aL7f�����If+*���Cy���&��vq{4絔�3lx�]�ȳ�����\s����F�
>��K�[9r�!u�j/�H���C�ħ�j�5�<O��ARt�.ds�������
��/�E�VG����7��q%Dg�6��N�`��T�����p��f�?���#
$�5ɸķ�+��������j�@�̚��32��
��V޽abIܝ4�Z�A$NŭĀzhZ�J7]�B�� ���})D�l��������}m���h�E�ͯ�1Q[�Z-�$����(�{�.4�P���Mɘ<q�D�w�M7G,���9Z>���&������>�3��A,�1�r6VOU��0Cx;��-o\*�K�&y��B�Iā|����`�9[8�s��=_|K��9��ă|x�)�`��X�A�n�����ܗ�.��Т�[��(K=֐ԑg�������l�]��cԂw�
�D�؆ �=1t���l��]KRW����I��nH����j��#pt��WR�	�-�
#�D��Tm�e��m|E�)\�E�L�S��ε���Z�9C��f�|$G�#]e�У��m�#�;�#���"����n�
�'����eP�6��/U���ӕ��;U��	�BN_�o"?�}Eh�_� ����J0Y�[�H�=l=�����go�t��)F���nw ��9ǻ\��\�"��2��P#����<Sb���n�X��\)�}��n� �k�����А�������/�ⷅ������0�D�@�iAy8X��͆y�1�������H��@2�c�p܆�7�u�:���1~ڛ'��z��|bC��w���r+��Dҋ��e!�Vƪ�+��R�*��U]f&�T�Z�2��rCT]7Q�j�m}ؐ�,3�"Č�m����|��u�7NlS>$1�\�5������ّ�=��V�Ɛ�*��O�s�\JQ����Qր�F����a{�Hp7)QLX͵�(�C�6B�O��CP���/z��	E>v��j�t�/ͧ=x��$�nv�ީ�D���Ls�U��i(ݛ����8�52�)��%�fW�b��Z��u�� ��~��?����� ���a������>�i�-�̓6��P�r�m@i�{��3�~����^���y&���&&m�A�ո�(�,��	i�	�{�h"y�L|���ź��DQ�V��f[h� ���j�GF>�Q9�y�j��[KN���=�7�)N���	�l���wEK](7����1K�C�-��?�u��C|I�|��Q5t\8�(
�y����	7N��0ʧ�p�.1y�^�lq��։bǓ�y{��*�p���������z�?�.��;��N��7�u��%9����\�0͜m<u��(���W��&qd��R���:z��W鎎'j'	)��������z桵��w1��\?�n�C	h5i@Aq�u"�S�N(xހ�?���9�I}����{W~�]��s�'���?&j��`coދv�[�Ye�.��W}B	����~�s�U?�^��P�(v�O���
�Z7�����SQ���Fw�#|%�k~��΄ LF ��Շ}�Ǚ�[N��h.��I �l��i]�,�D΋J���0�CS��{�ܸN0�`�'�{���_�r��9U4�|�W�Z�sA/��~~�==�����w0�����{�aEQ���_f:˾�.S���Z�\�Bv��/�B�Xn/��T�1���`͡�8q�u���2�Ds<�NZ�E�m4^��n�!&�t��t�&�!5c�]��Sk}�wW�R�N�ĕ�3*(0�^� ��������%W��X
���jf��2S���,���Z4�r�n=��%3�2���hA�A�R�q�-��d��0b�vx*�_�U�H
4~�}*L����6E��B(UH�Ǎ1�x@�tNႮ�]�F���oHs�Yn�C	p��l���HW�l�ΕG��P�=��@^y2�����Te�˰�Ǖ���4^��i�]}��%�0�¨��`�t^��'��{H�6��b�5V��bL���P
,�D�1~�ibh���9�.G1Q����<�	�q����%2�=�_8�M��h&c2�k�g�����>�H�'����	��y�B����P#�X̀!ƈ~��h�qy�*i6�U��kAnZ�'�I�b>����I%��,6HF�,Gٿ�s w�%/Rb'�!ބGYN�q",�[�ʘܺ�Jv�zn���t��N����̝�q�� ������1���h���\��4F\4���s��@�F͸a��ʤ�Z�_�0���Iwj����i����b���ǽ(�a���~=�����M=`�;�c��M�}���c�M�8%Ȫ�><ޛ�車��ʲ6ܝ�]\?�s(�|XN�_>���P��x�F����
��ս�K�%z-�ʹd��G��z\��.�W�$kVZ	vF�U�����c�]
T�;������?��d��+��a]s����\�\ƀ�;W����1�,�.�um��%M�6U���Ej����^���Q=���>q��P����W^�U�M���.��#�ٺu�݅�,�{e�%�D[m!'�k2,s�u��� �@c��8eG���-5ͷ�R=/y�?*Wu٥5H>�l������e�6 ۳��	�7hy46~U(���"e�Ec�W�'��L��;���bT��s���NP�'�݀ln�����,�l��jD����N�Y�|T9�eu�\� ��+��v*�m��F��i��fF�Kz���4C�_N&��u�_
.:uu�ZNU��ט��a��d��9��:aV>�`����zR�Wj`iA�E<��)�"ɂ���z^C ��?�w��b����o��A:e�H�p��}v^�}�-?��P�):�x����IJ15�KI��klA�O���zu@��J���������)�f�h�l~JR�ۯ�O)1�j��.ک�O�ȶ���=��v�#V���H2��@Oz}��?m�O��`��v��_%��_(�X�����3>��'�Pq�����ԩ�J`�{>����ON�I楻M�T��HԠ���B�U��H��@�����^��qP�����4~dJ@�7��&yg����A��UG���]���]΂{%��
ɼl����f~e����ݔ>�w�\&w�ő	���ұ�bI��_?��p�{@��q 4���r��S%��̦4�i>)uݘ�&rU���ւ�4������v�O��� �'�yu/���o�^F%����l�b�8�YR���EY�4��>^?J����FX�1����?0��X�˚[�(Y�o��J��uO�s�a
�}�a]lƖ�hA7~��M�OU��]Y�~��n�T�$뷩7���}$y���\	$U��E��O���e{�ً~�yvOB-�'^��}&�]g�n`���g[ts�
�
%�����a��I��^"��f�����>w���U�ʤ�ݬg#�9�U�[W�ۼ�Xm��G[��v���c�eFK9���T�Y����ճ�䝃�����M[��&�/�:Ѐ|��N2u2Z��#O��1b�_{5�����rz_��%b_n�?pFh�o�0�z<�$ȏ�R �����&�<c�An�#�����oW����&/�:oTp�7�p	.7;;�!' Iޟ�F�'k�r�bq
�v���z�)��1�行*DC�M��u7a���ax�A	��Y��9M����Efrٕ0��@���/� �̖w�l��7R#��rJ�X�<�NR�,K%�0PsbY�Z'"�����YU�Ҿ��
(�Ӕ����4*�6����'�w9Z��*;%��_�,��W�F4ܛ!��Xt�K}�=��՞V�h=�0n���zAI3c���̸�n,5ǂAG� ���`�y\T��D���)�8:U6t?�lLI���A�;�Ш�����s#L�s\�G��Z��2�'�i�c��R�������Q��<����g�im>k�`?�`��O|ڶ�`o�`s;���m0����_���$կc�?T�81�����5F���c$42=����`3�_�2��vHi���:�#�f0���'L��4{���m0�Q�$��Tf�/,&"R�d8�T��^iʀ��|���x��`w�^�c�]X��>}9�:�>�\]C�w�V~�=�>��!�5�\ѓ��iS��:���t<If�s�b���w�xU��.����>N��B<C��(���\5%Q�ܬ�3� aP�>��0���?y�k�0�f����B�Q�l|�!�|c��f�Py(���w{i�R𡗚�y%|�S�����wv�Gp�DQ{.9�}O�)�_�>W�����}��ea�q�	F}v�7��_s�r�M������m��A�9	+\_����T�͹鷂����!D7y`�;�F�Hx[ ӁU�5/�ǩ04J
e��w�(�pV�3U�$3h��hu�{@`��S�Jc^�W�d���a���M�7�R�:-
IC������W�8�A�D{�	��n����@�'%����l蕸�`(��kЯ@�|c:C�T���7-��7ӕaE�K��{�4��Pբ3���rl �Y��Zí/�O���,�;��-��f��^V$���1h�}�iH�L����&�m�2��7axg�K�V���B��c�S��v�4u���0����$���4;���><��8e��D�ն�/����an,w��A����i`���M�	 �x��v~�S�|B�`�/V�������X=@�6��PKXb&1�=:���]��e�_T>���*`�taٳ�%�7;ˁR�k��G�!�U��IX ͚$�d�v�d;[ k'��ɏ������J%vp��	�&���!\pX�[\1��2��-�ʂ+ :�p�A��7���E��$B�[^J��_7���~������)l��u�'�!>�\k!j#!]�
�f׿tM��@\�&U�yZ(�2j{��N�.lo%�I�?*�Yn!V` �K�{��Һ��ȡoe��1zU&T1ԧu^���F@� �>;vYc�`�N���q�LS�j�Z��  WD��?4�1?�T��9��X�C'���@?.ߡ�!�샻)�I�d���Z�|�/����[��n�$7�b~Я��)�ɘ�t�e��X8�M1��r�%��H8˂�z�)��g����h�SJ��v�SYJ�:�G�d��ퟯ[�>	�Rl�Ž��W~�"��]��Bj�x%�XL��k:�%����r;�j�A����E��V��*���o\n�t�`rQ��h��e���7�M�C�o�+�RQ��D�*�2��w�M
"�3�F���ad<~�a�YЧi�ފ˛؄������Z˕嫩㰃0��Ѹ�ŏ�%	ݤ7ۑ�����ob ���a�����1�}|��0�}��|7���%
�@G,fH}
�K�7h �0�|�\��{qzw��a���:� ��.`:(�?���L�]7@}���z��C�%EEZ���rq0�t7gǡ%�0��g���s#$3�Ɛm81k�0>"����^Q�=kEe��2΢HK�Ơ�L	r�l�<����@2 ��pX�� W�m##)��0!�=�+!��: �h0_X����ڷ�v�@�=�Oj�E�O.�2$0�=�V��m�[�H��K�o� �\��ݮ���0�����t�."qaY��>$�g
����G���SCRSNbjg��,h�e�f�~�Z��כ��\��A�q��Tv߂1rO���T�#D��j���n�_�~k��Ǥ��@(5E�[ݑeC�O��֙52ȷ��A6b���.*�%�w���{����:�R�R\ts��T�$t)�jP�9$�V�]7ڒ=�" �ԯ�1�{ �53"���@��}s���p�/�Η���0�r��P۰,T)�*�F�u��K��a����5���㻩~&�����:��im�S�X����B��c��mw9Ѻ�")��tX�����������:V�x��cݵ`7�nt������6�S�xDoD
#7̥� ��{�Ac/L�� ���i.9j�����:WR�+��������r�	����r�u]��//BT�pO�h9�4�IǄU/~�"+��|�����)|N�&�'�{��'�&)��YͨAO9�������ɤA_��GW_п�^�邥?��@�!ޫ>.�y����VgdѲ-�RzWZ��N}c���]X�&�#Lr��î��Kiyԣ���ݽ��PL9�JO� ���n��xJ�c��sb�	�v~Fx~���a�?ڵ��-�M��w_y�?)�7��,�
*�+~?f�f�*SHﻠPL7�\�{Ȅ�>��<�Go@���論�(��DM��w���`����ڬ���9B�>�Z�<@���)Xd���6W��)��,ɚ�u�,$����u�_��5����!/�hy#鉻p���P�5׼ݓ1Z���KCIJDT3��Q�G�I&�"	�-�S&�0��XP��Ý[DN��Y4ި��X^�R��K<���	�/}�Y܈nu���zHT�cl�YJ��@>�K��v*��֊�|���M�т���	7�%���Da>�O��v� A�b���bRV��K�����u����2�@�t���nBcj����9�1���9A�c��0]{ ��r�/y"�7�u��||t�(���|X���r!��Ņ�K����SRI!a��K(����Q���8~��.��8	�Q�d+(�N�P� ^��?�";�8����Q?�y3k;�R��aސ�ܸ���%�_���?ncT0���A��8�Bo��02�g�Q�U�Ok�����=�\����&���W�[!���$����xnr-��Y�Z��������o5*�	T�'$���fJW����x��a�,μ<��Z�aŧ�X���	�`����"��d��O�>��{_ʤh�52� ����L�r!���*,�D������bK[d6�.�uN����B��bn��Cٌ<������I�LR�׎ ��>��Rc�R�%X3/�0Wٽ{ZѧQ�s|�*�Y
��'�����RT]�&ġq^�㊭��-.,�����k��"9Ƃ++�4�?h��dG�7�ö�u��yQǺ��F��/BxЃ�=�����Y�d�;-$���,hl3%ޜ��	~��.�	�L�O4�'����u���w���ϱ�jv�ށ����q!���  �^�eI5�v�@�J!It�����E��t\`����(�^���`:[H�!i�^f7���m��
��g9�v��^]nYݹ���k[�/܍��S�$�2�4Vl	��j��Ea�-؄�_J��^�e!�)���o�$m�EX�Y,�Ǥ�Ia��#}��o.�H�R|Z�me�i�E��G��C��n�Sr1�{�a��A4�A�ۘ|��K_��UGL-��-�����	$>= �HZ�$p�H�[�`1�5�k�?���#N�?���P�,�{�C8ى7��-�?ď��m)*A�9�Ճ\+�*�0֑W+��-*�~�8|��$�aA�̷!�A�#����Vި��O�X����:��mK�)�vI��o�E<J��o���+�l�h�0�x8p���'gi9B�Ǥ�ˍ��Xp��������|yc}u҈�g��u��I'0����(��E�"]�_���F]�P'g��ZF.�9bc`�q��G5�M�1�И�46Y���� ��*z5u��y��y�'�z��U�=��QܵA�.�8�r��ъiC:�[�d��?�bNŚ�����f������� ?�à��*��lhވ��@�U��-��̳l��ÉZ���TbBoK�O{c5���QS�	���٘I<��?m��B�� a�U�/��Mғ�$����:XFj!��/���0t�Ǜ�B�ćW�<+���G�pm�1L�Ǡ"�y��5H�)�k��!U<�Dݺ#��N�0��:P��O��4�T����̭��` U��������Ԇ����x��z���1F@�Г1�y2��b�ŠQq���m~.��MVO!܎�m�}w��X2�x���4���4��R��m#�/��P��������y��N; 5ax��5�&��i����*NlY��Ů8A�l�k��vF�Ū�H�y���֏��̑��e5�ˏ|azѤ���P+�'�@w��Ū$o~Lؚ�0jy��AR^I�2.�T	k���{�?��i-s�������d�U��G<u�QMC�I���/�.Tۨ(�Ӽw����`�w�A�߆�
�]n�nX���'�����,&S��&h�ε�h��l@���D.�R�b����(D�kd};����.9�����M���Iz/`[@���g%Mt%ጪaND�Vx3�95��@��Lo��}ň��ё�'w��j���8:��B��`��}x�w�jr���$��X-V���xD�O�y՟N�g#�hH�d`����i
>s�]߳rA���A��	�7�ojΊ�2pxj��{�.�[��m���EY(�ʳÌ��~�Q�G�3�9�+�p��Hu�_G�l���'��ǰ����os�t5��
Ek�_���Z�o��彥H�����"������1�3� Lo����\��9$�=������/'Ȁ`�"��X$�:$g^��㋡̩��Mܾ�ee �.;(���R���9�m�� �s�]�n�*ZU[��:r���� � G���6'�s�xvT;��k������H_����4��R�lIN�����x�����4��4���LN��'9c���n����h��1�7f��\�H~*�N+=!�C�]�䣨Ba�w�t`� ��c���VǸ,;w��W`�u��V5�(��8�삩�2�ݷ�0����|�6[0�'�J-	!���>���>���]�?���y=æ57��\�P�tCrk�� \=���2@&JV�����u!�R��*��v}uAym�ᝇ��ȷ[���GT.����IH�/9i2.��~S%�T��S�k�|(��Z�N�pwΡ��eV�V�~e�	�pvx�tp�\<�
ȡ00�,���,�Wh>�u�1۔paGtfm�MʶU��j�����@rf����/3����#1_0o�։��}7�Tw>��*��M�P����A� #�C�=�.p�#`�d˅<`�0>x����7�\֕�>Z����l�w5�C=پ��Z1;����f��$�T 䜔@/�l��%'�(�+��ʙ�p�z�!�wv����Z��ொB�%t�Bi�8��I����4yd1����w�W�zt�$!��6��_��v$� �&���z����V�֏n�F�r2�I͚����R X��b��Y�Җ�����.��J2�ĺNE�p�d�Z�x�� �<�?k ���n����NA_U��)�P -� ;��4�xj1�=�^��l����U�+�G����� ?�5�"�֢�4[^}i�l��X[3HS�����~��5B}l��=}S�����A�����޻D���J��0/�a��F^=��ܡ�'�9ט2�c�2 ��ew��/��_$Dv���5 �kf��0���Xa��W�Im�x��5��i�Mj�Ft>� �C�d�v����$8Hi�ХV"���7ҁ�6rp���CRσ������D���7ک큵��0s��Z���\ZU{�	ۜ�) O���]Ww��Pa��vWF�Y�e������s�Y�[&I�&,�&�J.�
b�����;�xX�%|��2{}�ޫ�D�z�/�����d���A��b���� �����t1�¹{�+*dhúXn@!v�UL�.�N�Dbv�V<C9}�:��B���s�9����<�hR�v	a9}��5ZS~'D���s.|%GdʡQ���4ތs�|'��'>J>6h���;�頋ea cKj�^���I��l�]\�����8�<y���ܱ������L�<�؝�%y)נjlz�~>�<���W�IdF���<xP����C�Ḭ��
���Vb7��H��,r���Y���{o��&|�}�NA�T�K�!��?���G�8%���nN�`p��=*�Ru!��~9�	�);.J�J�lv��Q8�͵Y��(p�6�G0;�هhD�-��"e�j��
QcJ�S6��	q��;�B �/YŪNg2����zg�
PCĺg��ˍ����9͢�s,�K�D{5�U�{����>"�2�}TuZ;^�akeK�˾����C��Eֈ���5v���q�Kb�C���!�h"J룡�jN����� .�	 ��	R_�t��i�f�W2g "�Ӟ9B�!�/�;N�ǐߴg1��%�خ,��}���%��������g��ڐ#MI�9Wg����ї��O�i_�}1:�����)��i4�R^F��O�k_\F��:�V������K�����G^��I��)�j�����V
i��^�Q�3+�^ݥY���r�B�i��sʱ��G�Ax���_+�D�_#�:���U�	b6�,GN���9�P;D�\s֒ji�����p�i�沱�C��(��߽�US�O;c�0�*�����3Dï��^�FU�ٮ/�kw��|���3	���'���Y@�'\>��f}�b�]�����	*��?��E�\��Z۶�%�B����gkI%�i���7MRB�Η��Uw���j_�{9M�]E`n�1�DE�Q>��ܑ��V6�m��i#;D�/k�n�s�lHʫD�t㥨M\�5�wP[)�Ks	�I  �H��cs��(��.b,@ �s��a.�ќ��,s"� Y�`�Dʡ�0������5��@���JCs�k�gR�SԹ�<����j"�R�_�Wc�� �
�'�,�7y�H���vQ��Ӛ��;5&��G9�B�}5V6�n�^�V8��c\8�u�~P���l��#Ө���y�>`P�Zݎ�$p�	�����9�?m3*B��{$�a	�{�J�B�9�\��a���w-�(�Oka��}8��7` V���AK��BP���>ǔ�%��z��=|�f03q���e��a�ɱ�_׆ǯ����(�D+P�1JV^_�q[X�UK��c�'WoxFo���HRJ2��~�J(L���#I�l���"��P*���1�t��n�Fgp��$��*JC���^��tkI�v/��>-.�>ɂ����l�{'7Aw0bfVD�K�!+h앻�tw<��"o)��(�?b�����g��"#�s��W�*�v~�{��X'�J��IU�j��?�Hc�a,ܬ5�c罶 N�V��F�{�[D�������J��@W߈�o���(Z���_����}y����;Tl��Ք�K�D����`�C�YY�P�� ��U�{7��G2V���}� d������Y�uū_h��.�����c����¸�"�'nYy�Kg��~�2�m'�s*�A��o�;~FtӶ�iq�����i�Ԁuq#��l'�ۓ�5�B᫬�����c����`����kd�-4��9���a}D۞Z~��65Non�	*�`���?+��+q��	��W��iW�F���6H��݉�=����M]���[��%zm�xIWK@�����e�6���k+�i=M:�^�C鯒�`� �|�� z�|�f�U�$�p���Q��PEΉ����?y���$�v�M������ST�V�X���!�4����@�#O8���1z|y�+u�R�>�Gy]���R�kG��P��'d+AsM}f຤�ත��qOJ��ԅW>������e���̒���IƝ�Ӣ����LZ���l��U?�ⱌZ̎Ue��(6����&m���}�-Vn~��K�����(�G��tN�a�r���	U�..8��"�gW��~W~`@NQ��~�a�I�u�jP9���U�t.��o������m٢!���ssI����3JW6�������06;V�M�J� ���s@uz4i��������	5,�R��`0�Tybx���+8���sr� =���B��G
4ζ_���o��������a�`}я$��+��
b���{�N�I�+>�go�.�I�o̟�T'�5U�#�jK�b�x�n��wV�>1�����p����M��B钝�74��1+��ϖS�)��J��.�8�U� ��^T��K+k�U�X��g!�f5��cM��n�����T��n�Jَ���FV���h��F�ɦ>�[�Gk����i}��eJ����y�������C	��[�4c(!��c��W	�d�R�cI3m���Z��(��ϔ���
�=�kK8�+`��U�E����DDr6���K�w�������;�0���Z����D����,�x�̌:i��R#�E���vtt�
�R����k�#^qWo��]�͟S�;�0��z�(�+��~o��R�O5��T��?�w��(���c��8���ϝ �*�{�$F^⬋��B��j	�l٪R���0��4��1U���Y�K�L��! �@����L@�%$O=%��UU� ��F����N۫K��W�	���� �v��"��\y�S՟6���5(�wq&e�(�� �Vf�`��l�zs
-}��J{71�diT����ѡm0˽m`01�nMW��3�mO�K��\>&��%��b����&
7/2,@�g����LG�E�(7�� �wz��	����YL�=�'p��g� ~��gd:�������cƉm��^��N�lxF��z��۪V�Y\������|:��5��PC�sFd��{WM�)'��+O�TDhd���cVK�ÌBN�&������N��T���P�<ɨz�`.�@�@��ھ�AF$Gn)L},�'��E��*�z������.I���9� +��;�לչ���lG�#�R�翅���}w}�⯂� �j��3&�6���:4+X�&�mc5<��L��p��1p��]]��cE�Pi�G@�6(��(X��X�w�!/��`�0)��B\\��H�\Yܴ���a-V��Z��1�u)���3����D�]n����@�o^��:���d���@�����9���!"��ag��t�y�n�L���ɋ�}U9�G��%��O�T���~��{�.'s�m��ԏ�R�Ixj���]~��Z-���Fl��5�x"che8�|�X�b��:=��wӣ'� �+ɺ�w���D\4�UvY*�"���@-����v�V�/3t���K��Kb>���ҝ�E�ɬ�6/��q�N2S��W�|l�.?&� =X3)��OF6��W�x�}�>e��t�u_�xH)�?��HFg5{Gs���M1ÈZt;|9Х4yfc��ץ�>���%��Ŕ]s.,�6M�<i��ʯ����w�|:O��m.�Q�H;}T�J�B~���7\2C�k�d�i��4�t�J��Fh	H�UD���8q�	e�1�U�pwf_��x������*�愦1�bӏ�t������;�$�D{«���K-7j9�'Ð��J�~a�m�ѰE��K��<� 1�P13�a`Cn��)`�(�-T �ݜ���/pD�0�5�#��-��������&�zƈ��m��@��d�`�%_�@JMɇƆ�n�{P���\6�b�L��?�� �:F+-g�ˀ��a� 1���k�1�[�f@*���+�tu�:6�ia.���D{���QZ ��T^t�*�o��j��I#�Ϡ�K� ]��(ZS{9�Li�`�f�ҝnx�F�����3���4
;W��J�`Fv�l��͓4e�@5�,A���/���'���#��+�z�)Z,\vQ9���e�qھm��+�q�^K�����ÈP[*6��M(/b�ɸg%�ZU�nk��ē�������e_؋$S�������᜽�^���M��2�%vN�@"]\�}0%[~�'��ro�?{��	����cx���IEo��/Hj�mp���o��wO�p��) y��jM�ڮ rjrn��Y�3*�cb�\L4cӠ]�U��*-�'�_#�X���#���/��F
ꪇ����s`9�qУ���LN���,�x`�#[��nǺ�\܎wj>M��`�%��Gl���ф�)�~�%�� ��7Fv�\����֟�Bd��<��-;�3��2N�ۡ0w޶{ 2e1�DTU=�o��[hWѢ2`6GR���n��WYCzY��@�ߒ�>%�ԗ{�,kƒ�����4����)=�*����ֱ
n��>q�
Ti�<䭶	��tv�xJ�]�U"���A��;v�I���]Pn�g�"����~@��f�1�~�`�饑���l8�v��0c�q�~-/c� �=E�얋��WN�s	 (�~1�HF�O 2�dі�C����NN��K>Q����:GG��*烔z�-26�7�rWN��c��<���2($��ǰɼ�!̟�}�ɗ5�кU�WGհ������.�:�� ћ(�o�2�]��~G��b���CY����G�h�-�\���A J�2�z ���$0��iapM��̩	.��BQ ��懐��k���j�z�-��:�Ќ�:�?���y��q��ǆ��[�.o1�_��E	˓�'~B�r�k�Ce_f�&;&݇�#۲3�����
�.sl8��H?N�Bi��l'�ݟ�*�C��Ǹ$���?��{��\ڲ(~v��G�d35`���-�/g6~��s�!o�hT`�:�*�����I{x ��V �9ؙa��\�RTT��,>[S}��p�9(š��`�/Ơ	�Ra��3`��%�}�LM86�����5Z���
��2jWi���� 4eB�t��+�S���%)��(b�]��|�e�b#�
�\�໖'���&.  #��4���N�>��a9b��2n�����m�טq��|4-K�=����1�G�J(��5dV=CA�/,'��z\QP��OM���s}]��:>w�	�G��X���6�k�KI`m��}?���;yC��U�D돐��ݶ��N�@� �[�g�\�	g�G�7ZCD��D�3�' 3ੲ�l�����(7qe��[`�n�:�;2��.kS �A�;/������#$B�qo�b���㍪7�q��`S��Q����h�Չ:�5��LeQ��E���'r����z t*��� ��F^Wz�����	8�e:�\Њ��{:��Tb��rnI
�O��ã0C5e����;��6#�؟)������S���r����TCw��c���	p��q2��L��"�'�2�7K�q��G�C�_ni�Y����"y>m<+Tl�0�,"(����<�R���y T���(�l�1}B�bc����|o�0����,E��m��Kȵf�r�2F��������%`Fi�֔܊�n7�<;�e�'H3�U$�H�N���Ǳ1D	.���[���I�5�A�<Z���cI5�2��}���|%t.k�C��`��o�CMxY+z�ɟ�q�-� �7�S���ݺH�7�`TF��P���J;Dá$I��F*��b�cĤ�{@Tc�+hᴑ��l�δ{%F� )c���������=؅�u![7��C�j\�?���T��F	E�ߨ��(��1\����dR(š"������ y���	� ��P��Qj�W�iQ	'7���0�S|CX1��?����,e�ua��a�[���ئ�[T: E_�.�{H�����!j�kqr0��_���2�F�l<���/8!0�=VF���h������a2�i��e�[�E�1��\]v�q&B��d�k$��ldw��%5��F2~�������F���ͮ�.���C�W!�k��aH��I����勑�n�E��q`�톁e���YD��8G���Ke��4jJM>'w��#V	�,y3W*	W�pz�O2�����)2j8�a�Q�au�O9
�ܼ�f��
��9��ټ��&�dK\`�u��m���v�B����͐_Ɓ��YK����X5��L߯z@�l��)��ɬ������q��\� |D��X����
�'��?G:���&[_R��&�)�?��@R:Z��S
�(��h�<�y�[q��}桦s��o�k��w�|�t�ϩS�6���0�Z�V�*M�e�ߊ��� ��J���D���o��^J!�b���>̽X�u]3�1��-�陸�,Lݧ�gN������r�%�a���s�5w�%�:l) Vk08]d}O�������0*��*�{�m�f
y����]M�T�"��_]�"��^�W�N�E�Z?/�2=�9ߏ�!�O�n����Cj%��/�>@ �F jz_��39��ey��5-���<FjbF'��P�M9)<XXkX
Kv��G�²�����| ̎���e�Ȟ߹�^��"O�b�� �\��93��\ǲ�� ���D/*.D.���D�|�x��v7Tg�����My��K1~�_��B�9oI�=#y��bT��M(Ԛ�g�%�!��ʭ�Ӿ�93��r�#(�ee�YngY�[���Wj�<��}Щ�g�Z^iK��ɳ�/��7;��(�-���]�-����O�Q�����9�ԟ:r[:=����=�����Rs��
�D���x����	��w����`��_<G�W�e�W��ȯ=J��B���P ����[��~��bu�4ڮ�6���S��bsִ
�� 5�(BH�q���T Wک�M�R_�m�tSs��0��֨��s���	�c$�J�5����1qa���f��A��cƢ?].=j�z<1|4S��\�Lg9�Ț�Q���hV������ܬk�Sݹ،I#5�6��՜�G�ab�I<��N���,���Y���\�b?�#ģ��Rs��D�P���O���^۳^�����l��gR�k�������K#�;��(�qq�P'���'y��g������;��п��x|z�'��F��rJt�S���������a $ւ����i%^�b��"k22��5�DNan(VF�f�$�)���V��Oj.U��d?�z#����F�@��M<�Cvm=DF��3�����١�gպܐ�ļ�w��-���n��_*�����?U� zյ
}^�*w�/�S���.�� ������!�B9��Wߢ��7���i�?�q�F����')�cR}�����.=����7l�۷�s�}�/�Z�8`�)f�b�Ukb���M�p��������f��ֲG1\���o�n/\�7��I�h���S�� ���~�:�fcb�r^����w!�^�v�/�&'�0�i�t����fb��S�L��e~��|�<���{�9)����m$Sq�t(��d˚�����f�m�p��;�:5Dz�C�Xm[�eoU,�HV�=̧:P��9�{?�)5�2i-ʉ���.R���k�zM�� �2�[1)nǥ�&��`<A�͞�s�!�&�L��qp��j(n��  �D,�h�oJ�T�� >�A����k�V�A>����W���L�o7�j���q,����8&�h5�0��3�@�ّ�G΋X2ː��>�(�5*��OY����6��9�Z����; 	j�&Z�~��o\:{I ���TL���i>R9\���u^0���p���{�	���}�MIb�-=N�A�6��)�
�~|<C�2��?^|��b�b���B��口�svj�|&z'q͙�f�����>�z;�IYQ�|�b$����M	��N^���a
�״�����bL#R^�n�L�F�&�i�o���5���dY
�)j�A�ɿf�N#J��9M��^R�~RWi����4�5ʹ��&��
�
����:s_�5S��\ U1ю��i-������lay9����r#��Pw6]�!���������5"	�GӡA��.�,/��I̜/i7k�;{q���Dnmŝ�'�V�ן�G~�z��H�i�Oj﵁�*�<�]�A��%h�[�6��:���E����F?B��0�c\���u[����oeE�*Yd[�>ݵu�B���(��h�X�� Pô�M'&��qW:�uE#]�	$�\�ǈ�+�M@�k�'��� �Eׄ�p��o�S�����`���f�7O�����S�<�  bt,+��M��~S���y���B����S�ޢ�� �u���Dg�Vk�#�u�'KǮ��+fA�T��`���B����Ӟd���Z�os� %�����(V����	bU�"}_��N;�z}b�;��z��5���t.��v���W�2�?}9��*�-�A�(�H68���֣&a�ά�����-�i�O7'��'}~�Y�|�2�8�����'HP��q�-���h�W���������u^�N��(t�w>����8�-�TU�Eխ����
���Hն&������=/M�x�L�S>�~oN�"N_��d:��)�U*�ΓZE<��|�.H�����Y���%��T�k�kl����(���H�11������hdgs���إJ�P��k;��평O��|Ֆ|�:�-��<�jPz������u�>ܾ�D��Z��I�Ǿ�n�}������0�We���ɢ��"�������_��a?�����'���Y�Z�Cxc�"v���D:}`��~m^��<��
v�� b�����y��	7|�c@����+��#�Tn���[D��,Takt�g5�+��x(孋C�E�������T�Fgt�"k�Ο8���x|�H)��3��YY:��ei`�ʭ�8�ؿp�N��[m?��e�u�y��A�����)ƌ	9�nO^_&�s�`�Y���̩B������(Z�׉U�)�G���x�c�0�AX͂������n>��Cf'?��m#���>�! �Ɓ8wv^�ٙ1b^��?w�'���bC:����Q+^��~"[���qp^�.�>��P�w��^��!�Gu�����$� o��;�Z����_H_�s���~��R��8�-�i�xw6�wG*��yN�*�e��2th[mEwP���!CZq%�'�>������@s��/qC^��F�hE�/49q�F�sB�$}�a�(�
��Z�T����@���ǔ�h3xʇ~􊬅\��?�JWu�7=�غ�H�+S�����+}��(^�ii���$�j�U^���&7~
xr��e�'����R{-�Cu��vP�`A���+y8U.|*�6DI��?Ԛx3�k����-���Z-YzG�O��1*�F`q�C�72Dp�"�_y�]�9�����HHB�0F���� ���{$�66�sw����[O�݂G�4BX�w��6�ҝKM����^ �W��z������R p���Ð�{[Z�3���ޘ����*L�*�b*/�,*�K�
w����:C>���r�]?JUyl��t�@��c�J3�� G�L=�T>૬�d�ZC2���

6xD��g��Y���d5a(p�za~+$�&0�>��v�@n���u;k&���NTvs-Z����r�}	�P{���ż=u��l��KH���}LJ�\F?�������t�w<s���L䫅����F7�Z��D^�e�f���S�[�{�:7�������j�Lk���*ܿ��|/g��?�����
�6�8KL!��k����z�X'�1H���Q�N��%ώ*pT0��e����c�8��0��ʀ�d�в����n�䇦�ݲU�5ߓ��H ��������+�ک�v�4T�i����&0���U�j�� ����_�Q}Ց	��T۸!m�Oغ��B��h��|*�(��h���M��P�d�H�+�X�m �0�"/�)I��k���;39+!o:,�������Xk��:�:��c"�L������Rӧyf�~��ݮo r2��u����.�-��i�%��I��~k,���u0��v�j�+SA��,J���N-���'�)�Z�"
��Ac@��v�R*�*ievH>�A�T��!�b��}���I<ݸ~����L�9#�q="5]LܖYY��eW��������x�����g��`;��p���(h��^�VM]f@�;�]-p��̟�~"����kr���p&F�z����5��Y`o��[�?M�2�`8b?��Emv`A��j�o�fQ�@yi���)����g�x�iO�>dO���n>��ВI��@���7��Vެ�t ���K���	=�~ �စ���:H��i�և���e��>q����!ꖦK7�����ap7�Y�9�o�}J��:�K�:�E1��&�Vޗ/��7 �cdEa�bFQ.�����yI�逑_�ptu��6j��{2�&�����m���K�Nd茱���\懮���hR��8�����;1DOB*T��d(/�+.0��$�%�V�������:�*��@9X�(ڙ�]k��ώ_�`c�/eP\ X܅��+���}V����1�i�HnXa��8�d󻍣�Z� 8�f'D0���ǭ�1��8�LF1�L��X�,�
�1fl�q�B� v#���V�%�����[q���݁i�ԪD����ʣh�;�P�Tp9(�h�fD���*5��o���[d���%#����Z�B$�r�����u,<!��_���V(I%�X�M�ȕ�O⨤��Xeb����Mtp�S�A��[n{|Z<ܼ��Ɵ���K���_�֢�Km����ҳXS�u-`�!�cN�h����Ĕ'p4���v��K���wm$�l#����x35B�sE�r���q�Z�����.o�#J�jY���>��]�oI7���mo�TI�-��k��^�׃y��=I�*���S1cJץQ$9�9�S���__)��f+���t��;֗.Qm�H��ii����X�T��,����E6�+`�^wt��v_M�u)�&���p�5�a����;�_��#UռY�m��>�D�[%���Ú�fx��m(�(�^I�3�8���S-�g���j8(��l"��v�%�M36(U�d�ZzD��	��@p�1Ņp6`��	CG�!�?f�GF���;\�Fm��F[�;�D�#�ȭ�'3y���4�#�6%"������J�S��޺�M���뇈f���3�ڒ)�8�ֲ@Ҏ�賃��h�pFYw[PK�t�_������ÿV�u���@��\�Qî�ξ ��>H}2��"Qlq�)�d��?�w�����2چ�[V��9}7��|��M%��P�|����U���cio��*9a,�RTesE|�FYݵ�]���v��չ����f����O�²Ӊ�H;�5hm&��A	����I�0�,Kaj+G�H�f�i�ʯ�5�����e���s�3@���bv\��c,O��P�@�M0��f�Lr����"1� ��g�Z.��xO=�uz�Q����U��~:܄�w2HKg�p�d�A�d'y�Vo�D�u�3ˡ���!65��X�H�P�-�yrW)o�]�f��� �D
��xL�ކ��Z����%M>�5����l}ǲb1>+�z%޾Z@N��h��nt�	o�H��(fV��i0��p���)Rf
rI�����;��d� AࡷEc l6��;:�^�?kB��(MRI@Nܹ��|4h��v9��;������4#[C���#w�\��<��;!A�b{�S �>���I�ދ%����َ�#��%둈���9��2�4��S��>�X=f[ő�xA�<r*1}$ŏ{рY�T�-ZF(u�,�z:�/�8�=�;�h9c� r�j�h7��p�����r{� �p�>)>�LNM�e���\�ܛZ_1oS�+]�右Ƞ�i8��Z�$*o�^�4�ۇ�Ax� �>a��-#/E?fV'Ae�,@�R?�4��8��U_�J����o�>)`t���6�Q�6Y���2-��{��n�Y�%|�~U�J�j#��
�-C�K �������J-	�8���{5Ud�\N�*�
k���K�o0}������ ��Y�踦���L�_�~�j�8��'��G&9��S��=�u+�Ɲ�x�)9�:�Biyt}ڠ�����aS�_oӐfG��<t./�ĉ��=�o��<�^�΍ 0U�_Z7<*+��{#B��-g���x����Sw���U�TY+���'�s�3�HAG��n�<xڴ�WsZ��%��M�%�'���3'>��W+�p������j��a{ոF���F�K���!��o�#��d�i�<�o��HH������� ����ڏhA�M��4�߭�{�1��2�gȔ�|͝R b����6u����Sb�00ן���2�^G�gg��LՊ���_�
Ͽ�%��x��տ����.��J;_�}g.���Q+�:�(M���(�)�?�L,ʏ{,��u����s�N���ZY�T�k����"(��݌V��2Y�{�����=ݺ����M����ˡ�qS����.���gzU$`�����B�4 �(��n[�#��<��q�¿�[��u��^$$�<�}$��gm�cSc&+ײff��&��E���S�cB҂_V����!��0�I��J�I��wZݬO�	0b�.<t����M��V����6�ߛ���Yc��3��.K�/��q�T�ܓSG?�_2ts;�h�������=j�8!���n�L�f��"�����3� �S��/A���yS�E���L�{���*�(a�5*JԒAN��ڿ.�Q��2Go>/&t�C�L��g��k�h���i,�W�(�-D�,! g����b�j%�H~�}�_��~]2J���L�2�°���}В��b_T.2z�a�s 9���$������i�ْ�����5���Ԙ�g�Pz���=�va��ڞ����y���8���QD���Yu�'A۪[�}����7nn.�IH�G��SV�th�i����I�U���z������D�˘��&1���<5�cŐV�ǿ��P�.��4�ɰ��I�w�,_����n�5ǱT �iv��D69) U �����QQN�6dƽ��w5z[���O���XEX��Z0h�P2D6/f~�H����+�:�G�m��A��ͦ��Ok�J��V��J��͑�������e�9X}b�'{=���7dV��G��CshVH�ۋ�.h���j���3��gqJ<)~姝��0�wN=�}o,z�sbf�T+�W���.�a��6��@�����u�')�4K���ru��{�7+(�4T�+�4�A �M�UX�
D��=;H��M���0z���vG<`?���5��*87�ϒ0�+*�tu���W"%�5�u�lYo�l80�^���N�`N��r��pi���V{Z�M8�R~��%�+�.�3G��K�8}�`c�d�!z�9.�4���1���IGw��t��$����cVx�y]�=�����1�.g���9t��^Nd"<�2�˓N/�������vW|���vą�Y��=�����Ba�Y,U�vp�;��#�~�����d�"�� oV��*+}�b�������g�E= ��c�o3�eF2��$a(8���&;�0�|z�\<L'<�L����:S�&��-�N5�Ek���#$j�Fys���g�������bHum1ts
b���ߊ-ǂ[D
�;m����_�����=��B�����0h3�'���+�|ƴ�_J�Xz�L(J�С��j�u_��8��ha`��jl�B3xT��H�|�|�xA�%��?�7@ �!B^?n$���x�o�c�1�?V�wG]1y�)bl9��B�֦��񯾱��t�"Cqn^r[����1;�=�o"�6�E�6b�O)а�Ai��IiC��r�Lc� ��9,��i*qy̸e�J�VjB���Md�箻�&��r�P,3�p��Q���^���	�,�V�z��+CXp|S����Y,�����DH������E~�PEL!/�7^�4 �>����
�3�jNѝe����A%�J�n��s�Nҥ��rЄ��3#RF��&GLlU�~��f"���7l�5�Q,6ׇWEF�os9������fI�>N!]���Þ��2��zuO0�KX����E��	r.%>���~F�7�q�z�(�s�~�������
���a�{[�X�$�ޝ��-�!J��v���h[m�[�˴���**�� #���t�5)����@��6������)G��K�@�GjWy���4�LQB3E3TA�m�Wc_#�jʋh ��P�_�/����T��1�������luq�������L��%r0�Zb�����t��Z�:��߀��B�?�Ű<.BX�@�<_�F �Z�O���T8�(ܵ��bQÀCV�1�ɲGC�S���ޢ��?���/=}��!�
SG�&W�����ݲ����V�nt���$�II����w�!�E�U(�
q�H���XZ����s�z`���S����r��a;�V��3��˥���uވ�W`Ư���:�eѤ��FZ������v1���ٺ� ��󲆺��]���nvN�b�<�H�'�TŮ2�F����3j��֚u� �؟ډ? R�]��X��|���eJN⬑_H 0��Z[��MiwN�rδdJ�j�1Y~_a�8؃CO�g�����E�����UU�0i5_c
��;�ⷷ�W=�NF�2������zh�w%�?blc!)W)>�#h'js�~���J����W��d�4��M+a���`���'b�g,?&] gF:<�4Y��N� {l���2
l�AhP#�W~�u��z�/83��n�F��J��qIC�~���Tl�)�����m��Xx����H����EW�*�Q����ND�n�F���3#1�M�0dڣ�t�\����Y-��Wq�W����i���A��6zP界*3�=Smw*n�
��+@�2R��WڃG�b#d-�0�agNA�V������oJ��X�԰��y��uXu��t�l7��?ˉ�K��h*�{�fo���\$V����V��C������)Z�O�S_+?h ��g�NO�0*~� �(�����l�u��l�U��	�IQ�O[0����q��<�6�!L�7v�x�ۭ�{֪��)�ΰ��c<�tz�6T��XG�p]�u5�f|a�=b�Z`�l���Km ����і��J����{� �nj>���8�KOC�Q�n�>qxk+�ğ��������~F+�BH~Fl�ɥ������=����jJ���С�f��WЩ͢~���/4*�:f\d��Z��i6��9��u�a�_��� Ɉ�º,�u&�����L�G�
��{���L*���R`�̘����0+cÙ��'Uc�I���W�x�[g�84���g�D��V��w��4���ر���z�9��;�ow�����:����I�=��E�"ߘ�]������g<�ys2������%�S
t����i��]>����>`�_rH�ر�m��� c��`^�R	�S��j��!�����ߢz�|*�$��8r`��oL�|�X먝��I��i���e�M����ޑ����d�A�)J�3�{�O�XLX��.�؝�zD�wO�HJM�'��t"%�?�Y�]g_e�@�XP�g��,8�qg��uDr���qA/����������;�Q��<�ı{T���qlF�̓j����y�"����$����h>\����]�J���7�{�H�L,��~3R�8�Q�t�]�q"�/��FgkZ�bw�C:�����WY��u��+Jܥ���t{�M�ȃ�.�gt�Zq�^z��~�ٝ���d����D��3����$2Q�Y	n�un�����V��/�xJ�<��Iʂ�J�T[�A ޷��SLA-$�1.�I Q��oD�w{�l�Yvh)��]9��	����t�-���S��3P�$��� �+4OΆ�`�h7,Z7=�w�_�(&GQ��l0�;<}�kO#.��	 �{+�N�Zt/
�
e���#9�,\Y:uQ>�6*p�8?����_��o��?��(N�$Sf<EC��~n�w\����8,�e��Ŀ&��P)06�׀��d�����M�w��H�����>���Z�E��u������#h�]2�ohi0�p"�M��X�[�K�����2Îp�v�1?Y� @p1Ar�5����zS��%A���`<��kT��x.䠤�n B��(� ]J�_��#k�wQ[�;:�e��3$����������H?�Ƚ��I��������y������
��Z,, -���ʟ׸��k����r�Ya�]}:I�P/u�kzk�ԝP�T���g��l����j��J�T��t��4��$;�лC��O�i
=%t��f��Y�ՙ�H��x�j��B4�F�b�\Zl�-�������Kɵ��t�)#[��ڣm�j�>�f�7X1�qF�W!�y/!}�QmyDz��_�ެ��ݧ[�*W�m�=y\�p�uII��x������S<���{����d!E����+Ǘ�\I��3|5���X�a�!���%{��rθ����\�Y��� R����;��iA�k𦺬�D�/�@���A��t�g�VF�m�01��i��m)!�b��D/1���b7��;,�"�b5ڨ�*�(=ae3B{����x�.�����Iu�z �����3Є�� 'U��ܬ%���c�[e�ף�t{\�h2�%kY���u|��
rP9r�u�벮�������\/�"�&�1��.G/C8Z�4�E� o~��ɹ���?�'�V�j��UA-t���L�;װ4��:�y˔*�ea;k�k ���Oj��IOc%��p�q?vKš�%Y��$.wZ��W0޻���4}��L�=���P����&G�4�$2����p,�lc���s%Ұfj�=#�	F�~εc��
�M���Ą
Т�TA�e��?[5��NUtQF���]���ARt�1�ޱ�O$wuɊ�j�P0�rL�$��D���&}��%^6�8�?�Vr�I��`\��%�y6���Q�j�:k����о�TQ�R`%�a��8&���6_����l�~������<O@G];d��%xo���$�������d��	��A-���8h�~��~󉐲��St�U��;������-�]�u�&*c�F ����-W�3�	�zFsUs�.%{QF���6�g"��#�^��1�y�|	zX�����j�(4m�B�j�$LP�Wp��C ��5=�W�TH_������MB���P�������5��1DV�~�A��+P0ӖQLo��<(��l��;�Ѿ�=9b]Qv�My���)7R�����׊@�8���:�8�<����ˬ,G9V^ ?�NE��������$�i�O��/M�Ro*���o$����'d�'�|�qY`�QQ�>�����6�"�����"_���X��KTA8��H�f�Ui$:U�A��\�Z����9	�$��_��F=�&ԟ "����ޖ�k�����Ĕ��P�{����rUκf�+��{nϕL�F+O,I�UJ�Y�5=���a����-�k3c*���ݣgWF�ؑ,�y���0b����8����g����/��9�צ-e:;���d4��PP���V5���%���A���Jݮ�P}{͵b	j�C[�{�w�U�p';�ڈ�瞔[�����a>����q�����c&�f;�������0,A�t�bB!��#���l���z0��>;�o��� ��<\����[\_��J1s�B��G¦��]��?�g�����!�J���:g^��|/��/��y0��-��Z��~\鍊5AJ1e{2���J��r_�� #�sN��nV#���VQ`5��w�	���]�wE�H<��*�q��x36��]��qL���\-#��*�'�|�]ޛ4�#�m3b��e.Z�bG��NȓYd�e�԰A[���9]��Q����$���|��@�g���iX���ο��$�Ћ�i�1�fBo�@o�"�YL@��`j�N�6˱��y)K;����c�i�@@U��b��0U��y4�n8:5�ʓ|��"K����2�6uk�ޭB���m\�C�7K�f������h�6��#��ꀢÁ�m�
����ү�G�KG�Р����3�&e`�?&*� X=�|��W�6s�]�p��O�W�y����/ �f��/���!�0?q/.����vtsEt̻�+�Z�.Z���rd8���d<��(Uj�^���#U��DT?�p��U�`�%�$����̔;����%C�]b�o^�8��@�΍��b��K;*����V�qC�gM;����.Y;v�0�Ȫ< ��Q��!�����&�YcX���BN�'�����J й�� �!��1�|��+P f�Y�s@�ɘToG,ݘ�� ��͊���E{�hf�1��1؎�֢PN��fz�L�^u�����Q�
ztΕ��G3��徍L�O�H)�p����i�ᝃW�3(�̎��F�ѮDj��&����l~��\�R	�A4��I5�7{B ���� �,�[�><��q}���_m��/�5D~�&2Zg��R �tZ7�H9ew���SxVGURw�i~ǥL���R�S��� ���0����l�E�E���^f0A`��P�7ᇑ��y�a\
SUC�Ա�sOP�/v3��,IN5��A�a��-Fyys3@�TX򱢄Ku,��\%1�1ji&
�K��������,�
���zy_2�CsH���e|F$�&t3�R�������+��fp���UC{)�`��]SF��w_��y�e�k�G�;�65y*�P{�:�2��L����|f<�>�[�k�	���I�:�ՍH�t��i��O$��� ��ާ�H�W�[:O�hc�q��ks`2Ҥ]��L 6Ta��FY��0�)����.G�J��a�2�[|����1whd��/����<|���f��Q�CƊ?�n,�}G<9�K�T��ջLB��t�ۛ��Ge�3��������,""�úv�Fx7e��P�H����|Ą��CO_�'X�3#B�/+\�ȋDeEɣp��9_$[�uS	�S��t�9�ݵ��a3�o���`�M�H���w+L*ۭq�4W3{�͋�Y��KIz͏���^��7��lw'�5���X0?��Rr���<?�'��?�;M���ִؙ�M'��D;�
ۜ4W�E�%R�* ����w"��y�Zͩ��7pD�@¯z�jr'S��>�7�Mo�К�o���(>z����� �t�6I�Ts����E�[#���2%�d�˃��u� ���a��r;=���?�`��D��!�X��l��À��+��V����Za&3�5�IЩ/T���(�v��|�	�
�����W�����փ�������d֨ph����
��w?G�%�A^`�Y�+{:���e����Ҥ;��m�g���ƍ�k��Χ�"|��b0� �?�ht3R�y�U��CP��nj3��V��Pt���`H
��*�ױ��MuiU��`ڿ�<C6n���� Z�?BZ��GC:¯��Mx��E��m���fh��r����xn- J��@�Q �ͯҟ� V�4N��Q���v�������@�܋��n��栘�Du���}��Y��������{���E�2���
�$-#▁�2�F@��Y�	� ��.m�x<�A�W��/h�n�e�Q��T|fٽL��ϯ7�q��3�G:sv��L�j�,.8Ă�G�x�#�1Q<�kO��ǡ����L�SR�E���S>�l�/Y���) ];k�B	U��"�Hp�~�\����8����U<`�	,@���\��?�j�^�hv���q�:yŮQ�ƽ��>�e�.|A��y� s�l1�&��#�*@�5l��p���,��?�j�A2x�Ik��6�^��Td��7�����|6^z���;' ��w�1�̥��֖��MI�5:�#D��Ps��2�wæVʑ[��t��њG��f7���Yqѽ د$�A$����2�	Ԍ�fCOф*3O�:w��
ō�~��\�=(��)97��4�%$:���JyxY���Xw���xh"�jW<��c�q�2Շ�����;0cF�؀��j=�!�@9 ���K?����z�U�������poou��n9�����ו,r9��5�|#���RcQ�P$�7$~S���\UV� W�SR�0�`\�)�7K��P��pĠ�h$"N%�C��X���{���\Ye� ��x�I4vX��_��3���O�����9�D�!�<%�GI��D��#��V��]�{��_o��cl�-�kch?s�L4��y�F��&[J�_��@����:���XO�N,�&�� ���U��P�ej&n"E,�.k����G6(��<�2�\cF�tVEl�-��&^����f�5]���+����Z ^��q{�>Jl��AT���}I��k���y�p-�/���E�l~
D�kJC�q�F�x@,t�@��YW�D@}�'?�YF��jO%�d`���Q�k������qO`� �jsM4�m�u�d ��^�f��Tܡ�Bђ$�S6�/���!ؾ�>�5v�hʺM!Ǟ���8;ۣ�P�8����΢��F�?pD�T��÷dc_]re	�v�9��oGe#W�c̯waF��|���"�!��C��8�N��Be���R� -��NqikI�+�G A��=`���U�-�ޔ���D�v2+�,�D�h���;s�q��������#�򨥾$	*=E)��:d-2��zF��*s�W𘟶T�'���m]���CU}�*g�Ik��!��%��]!��b�yTx�xԦK\����x�\#�6�������/�J~ 1�G��}	��`7c�^�qC�����w$�z%*�Y��i6k޴f�D��m��%�� ����d�%�1]��%羽2�������s�	�_`�Y�C�:4�:�8��39K����閛Ε4K�	�e��q��y#�v�0p��29y����\z1�(߻q�g�U�&�䵵�Eb4 xO�D��.'J���S:VkQ�Ƀs		�/3NQ�?�O�6��;�	�:⺑;�T���s"*kgmd|��C5�m2�Zw3����o��Y�:=�KղFY/�;�_�U�nc��h(d.�Y��=�I�l��x��Z�	�];e�f*��n�t��s��/�1"{;�2����>)HI��
�`���$�	+^�W��n��w�Uv>B��}���0{�3�|G�%�/�ǅ3�[�6��L<	�3ug	��}���q��0��R!ȗ�<��XSvV[gA"����b�UBAȮrmĠ�1��ջ徲�-��`�t�Z�.�����hB'ȏ��cL|�|��'�4���j�y�p&��'�	�G�d���ɪ�5 ��!�X�R��9K�����g������#ŗN��j�H�TԞ�(�֡��O/�x1��a��^��'�-x�j	:�7oΑ��vv	�R��w���V3�O��t>I<y�-��Μ%��ytX���W���Y����a�y��(
��kd�TO�|���&]���,_pߕ��~T��Șk#ɉQn�)�v��Z��Q҅�g�k�7����WO,ш��oy ���d�^<R5P��fw�2�>g�j��e�?B�G[ _��B��g;O ��~����l�s �б����Cbr���:y%R�����cq�;��Ȗ��ͣ�����څ�� ��D����E��.<���l ��A_�&�t-��o9h�(��Ȏ���E��|�w_g�����&��z�������Z@�'�LgC��߸�B2���A	���u���"�):���&����d���5����s������d^Nv2����/��]C��&�	1G�/��o(O�c������H�#�͎Ҷ*�d��J�m��^�O3B.����#/A��u1��b��i�(��|��N���m�7�/�_����T ��U��k����+)H�_�%�G�����QO���`j<y�Hs����B�c_"�)����/䔼�8ӍZc�j�A5 �4��vX/x��FW:O3�2�g`�YTmlBZ�o
p��^��@��E6͒��R��Z3<!"�$��L��C�?�/v���+�� �i��V�׬L�|��_f���i��pR�;PH(��e��G���n���^�t���|x�zP��?��$���V�\����$ci)�6�=*KOx
:.W}���
w�}�/xsn�4
U���ڼR��^s4O)���f�&�y��*�N��k{�ڱS�p/(!�m�s��_�8�b$`��f�MK�d�w.lf.�O��St�^�y��vSU���N��A�ϐ$��#0��g#4��^�������ꙏ1��������A�';�;�v�úI>�H�Q*޲��7��ӑq�ᦣ.�)J��k"�xn>�k�����&���nSԶ/W���?{��kQ1�-�~?]W�����Z[���و�zܹRr��?E��n���0��{_�����ya4�:�u]8�`V=�%�g����%XK�m��2�K�k���۲�PyJ�0���+q��x��T����AF�e!�Y��QgU��rO�Sg�e��-M""����wǹ`����3YR�%GEj@��j�����G��@���N<�G�L�B�&�逸�O�3q������F�@�H}H֓��z�U��3�~C�S�����!	_�VƋ��cx�e�Z����A�`���P�!������ ���
�{��o��:��\=���-�!7\.-������B��	�|�"}��F~mO`��{D�tw���������o,@ �JW�:�@a�����o >�t�/K^	���U:�b���.�*t7�-N������2�FN���Ww[s�>��<	�CfX|��f;��r�[K�.`K�������� ����4�Y���TnͲ��ĿC<� �92�K�	��R�s1����$�̵�V���.�x�{m�!��\|ᵕ�Q��� .}d๬s+@�h�U���Y%�����Q���G����������?��"��z�����5��s�8���Z����7�U��e���+wq�o�*�T�󌐳��`K�(��r�b��G~�sDaW���8u2Ȃ@3�1י��w/"o�=ue:��%���� O]�̇X���6��d-:E��0Nc��؝�'���_�rގ�1����gO�?@s\�;S�6	JTv>��J�W�L �v֤������t�^�OCL�j�YL�_�Q\Z�tB?cOS�upi�ఴ�����ܰ�dG��H�$���M@�P��F�(h��*z��{�pIv����*�r�����|����sBh�/�������`�nVYj1��|>�3?]$���T����u{ч�Ұ�R�Kn�Qx�����kK��o�{v�l�+�0!#c)�E��f�?�L98�%�V_��V��<�q��Nh���m��� ���J��W���ĺ=+��<��yk��b�4+�J�2[�B=/��t�E�]�n'������+�R�s��6�7�A�]���ܦh.퐈#W�gD3G��E����)vk9����+2��u�l��E֪�����H]�V��bM�n��n�Q���Ψ�U�sB� {_0
�E��V��]��C�C�W�'Q�#�\�Ӥn�	kEc�\>��[�L�!Ryč{�%�R N\˦��`"��HZ	��I�>�G�29c��"�o9�l�����\10�ThUF_ɅQ����n��~��B�Ŕ��
DTk&��@��ï�<��'���$<umQ�wJ����`ҩ�p0�Q���<@�2����z�Յ]�����y�&`��W�^=~��A͂��$���*2����͛�3���c�}���4��5�~3�'�w�����/]��O�R0�S��k�M��SBE?C�3�#����	D���J�S띚ٔ��a���z]���ǾēhdR:Ŭ����TGn��]x+�#=G����#+>u��g/�c��U�D��s^]���ϥHP��e�����c����u�~zܭ5�fg�"���݂k�㪞�����w\{K�?�%mH���@QqmB�Kp0R�+�IOe�A���貭n�Y��_��
Hz"���v�]}��p��i�i���7;X#�K��v��n��P��.�V`� ��c
��	W���d3I����C�>?C�pj'��Y��怜J��dh�q�&�.�� s�50䝜uU_�Iy���G�d�pn�|��c�7eb$�*ޡ�/�#X����԰Y)4���(��>y���r
U~È�ë'� ;T��m��Đ�a���>��	f�kU�F��vJ��Y�uË�`oձ�*c�����<I�u���xU	��xl��I���&����`�1�js;�)2d�����������Z~/��Q�H���ȴ�f޽��u�����뾷�ζTA�6*٫ʥ���t- ����H�!�K ':�s���N�����H��#�HNMX��|E�e��H���7�8
�����WO0)ᶄsHoҙ�w f  �"�/X��1�:�T��'�&�������Y[��D��@������ʼ��C�w|��z�=X�x���N���i���;^�P���1���J(!X�㰝:��!_�d�"�'ž��d�0�%� 0���R�u*�*�1�4�ү��E��*��ڸ�6b���^~P��K���[�m�:�J'~G=�}���Ȩ#��r��ώ���X�=�]m�P1q�㌦���&�0f�&I3A���sZo)-��J{ =������&I��C|2}�����O��v0,C�� fÍf;���������T�dR�>򸥥�|�'[�2��p��1�6�VYxr ۔̇�^
�|��8�uOh�P�3/k��|]��51}Ȇ�zd)%5��#�<���U��ߡ@�;8t�� ��{u13N��Fˋx���`������Q�'�L&*-x(z
P���4a���L6��{1���?tc�����蝉�͕t͍d��Oڢ��T�oCX)z��aC��h�ه�d#���TA�[X���d�Z;V�I{[4��3T��w��W~Y|H-�<���,}ݚ�Ke�#�:r��D���{K�48		-K�0��4�#�>�Y� ��aRwt�gV�Q5���/�
o@�<�X2�z���ٽ����W�&�Њ�=�N]��!qZE�ܮa�=�Gۜ�x�j��D�m}�q�\�a�5�ᴰ��&f*D��V�}\�.p����8�z�]��P�$	P��gz\3,5���z��*K�Md�����~fE�F��յ��і���58���v��V���WD�}�/c�ƕ�  �r��������b������t'�բ�9'Sܐ+��S�F���D��a<���d���j��f�G0#�$lX`D���]Ow�U�lb����W���?��M��d`���h��gq��2(�qW��=�*p;�N��Y),U��Z����᠚�ޞu<f;~�b|�*V�'��n��g�"��ѕyu��k�cUXU	��d�b���J��{z��l�����
2:hվG���\��^fK�9ѻ���C�E�9���K�����rϬ��=�x�������bP =͞�Ӈ��C�	�d`̭k�E3�`ڑt��9�F��+l;�ץ&h?Lv����}����=���cv�N7�H�$�+~�m�L[�q�l��k���ʪk*U�u������y[66�mb�?m��3m��P=Q�J5��R��?��Z�ݳ�J�_�!\�͙UёR�o��5C,P׭��ƎJ���ew�hd9�8[Ώ�ݖ�AN�p�Ҡ�:�n&H��F�*,�3{v�o�����@
lG�q�_�Z��-�e-*-��;����S���k� �n�hc��kx��E{a��}���F�{_M-M�;�Jw��yQTXv�����&�ih26_���q�vy�� H^@C�@t��X3���S��>8й��av*{Z�e�2L��G?k;�XD��ٝRku�t��l�E�pUaǩ{��ʼ��=?3��F �� p֩:*������##���F3[�V�'�m L�]�Y��WR֡�<�d�n��L�R��@�e�MA"�4c��w�(m�k&G��z3B�Ď��{+�,Rvst�{|�5�3�!RS��@	љ��tؗ����d|�����8k���سi}tí��4Hڈ���d?�?	F=��=�B�Cb﯃��-7-�-:tE���˙�T`/�@�!"��G�!�!��J��E=����m֣@����@��"�<e�
��o���=�_F�������^����=2�����U}t�����si���/���B����#/�����Rk~:TH��qD�>|��f|+K,��y���n�����$^��I^��Cǒ����Y���F oS=���;5��k��S�[^�C2f��p ��]��F��>�@��5�	F���?�d�=Q�=�y(=-_�b�	N��n�sY�U9�7o��5���#'��>�߸��؃��,1�e#o�,^���U�^�%��V��?�@fZ+�~C�ל�D-���`8��v)}¸�n	����J7(� _~!��<��Z�yw������ZʰWBLWzu���V��BгJ�ⴵ�����Ri>�iM��b�j��h�z~W�=�Liz�>�j�i��Cj01~�vj��f� ���D
0�j�����@�����U8(���g�d��'ɩ
/7�i�=��r�w�2�Q?� �K&�RZ����l?�Wd���E���DT�rbH�J	(칉�*��m1��Ƅ(����16��J���`j�B�,�q���E��Az�b����C��U��yd�{����L�O�č��@V?љ�H���@ŵ�Ĝ�_�,}5T���¨ܝ�F�RL�D��w���)Dzw��0U�ņ�
�&h�r+�s�0t�9":�@`��=t�\��8�����U�2�}�{�����9��d��D}AB6�ãc�/�n�3�Q KN���:@|�v�FG7!��J<8�W=K%Mc7Ё∱��b���">/�4K!��x��U�Ϝ��l�"�xT0N0�k�=H���qƏַ~�v5���4�xkԻf�2�Hܧui� �4M������2%R��bN��._	_�"���xx�mQ����`��[�P_AY�8Z�NW�,��F�,;� ۚ�:���.�a,���E��U{5��H���fp�|ϙ��� �7��`��^Ac@ �)��4N�c�KV��ƭw)�`)z5sB���%�4R�BՃA�Eiؑ׊���l}/��9B�[��������aB�eU�}7"�#��9�:�i4�/g�PLH���ީ����f����d#6Aq��ٺ����$X4f�\SX&+��5:^/�M�� ��zw|Y8��z���x�(�����U��P�ۑ��+����Z�.�og,�%��7/ѫ*XB����$���^6��c�����f;A")t-`���CO �j-%�4;�#����~���'р�Z�a�/��ښ�M�G��ʅ/ߊ�ΐ�)[񀠑�Mۻ�L����Z��Xnڄ�)hx0�A{����d��[uz$9M�^j�u?�����P��61[�c�+��'ޣ��g�3���o��}V]�Ai�)�����ec}�%���u�	�S�Ln���`TE�/+�l�Fg�b�0ɇ�{�*Z��;-3X�|C5������`j�!U|
[<�6�jme:SC���,;[w���e=�ǅ5,Yn�L�V{G�����E~)�B�U�>��]3�"��JZ�v���{��1���,�+6�-���2t�U�pʴ�U	N������p�f�
O���פ�V,;�\�P+�d�?S+O#�q�3J�}�cH6���QSÖ�V�\���._+�TIl�r�Dz'�!�!�S4Y�Y]�uj�W!7D`�jfeLp���*��������i�u�>�����uF���������h���kֽ�Pyy����m�_J��.�>I�V��㑂L L��"C��y���0�O�W��m�bh͇up|���A�t�1̀�Un���	�&zpH�I7��]��n��)�;9��� `���i3���K�-�~?ť���=��,ks� ���7�"�YO���u-��=�"����wE��y�g®V=W�34�]7�c��yދ� ���?��*	*��~/&}q�0Cz�^L9�|o�jUx�#W���­�G�.����,�B#�a�O���T�~.��//�|�o� ��aF����w7��ktC3;�j��Ľ�;8q���2d����g�	nH��zvW-��%#�8U���ө���U���&�	�2�ͳ�Y��Nn�u)X�X�C�T��6kI����ͩ.�e���l�P��En�&2�z�x�+6��Y0����_����4n�2���i�oN��RΓ� �gK駭w���	��^�iD5�M��u���C��X���ԁ��"�|Σ8�k�,7����d�
T�η�q�?ZL�����?�N��0�6�4��!���lK��Z�uobL�#�Ս���i,c �F��������������b�ʹ���E�w���"�~������ �F!Ԉ�����13�<���/@ם��0����i�"A��D.\'��:�N-*3㲷���,�1��Gd�X��:�h�ū?-M.͒&ݚQD���s{v���D����z|ŏ^�P���9���.6�ЂR�❃�D�.D�B�:78We�[�Z�!"&�!"�]�.�����t�����\�0���=
�Dj1b�����O����<�D���̊d�DwI����u��8����K��fe�%B����?_B�x��������E�W_�!����A����He�qV�(9����4�Mz��G�X����M��A�Q��H�z�
�X�'i7���� ����ش�M�&y�w��)ݨ�Ҧ��!zr�W���;��Ÿ#��>�הF�"��e�1�����R_ߗ#����/&u�^	:�[Ny9-�N��vFg��}�ŭ.��� ��6�o	k�k��z)��e�z�yL4V�CL&H���}�ιn����a}�{�̬�{�0n�7T!@����V��O�����@jc;_��#�i{�zLa/��E�`�=~�5�5�ꄃ030�"���6�<<������'a�,(M�j��.t����� �D�^���땾��P��������^�����ر��X4˼e~�i��,�
�@N�yg����tڂz�MڶpS���i�9�>J'���_�!⨛�]��1{���~��~��q��SC�4[���*evR){38��x�E���0�_�����=�86ѳ�WUK��38E[�u�՜�g_$)Vl�M��e ��R�i�#8}俒Eg�E(�cE>���K�#��3F���}������|1���t|�X{��ϸbɮX�|7~�A�T� �%X�H�Ӧfq�)�DX�s��r
~ ]�}���(%:�zŜ�6�?�Z-��f��с�I����u��R���w:���Sv���¼.���-�Q<_�=�i�J�ηTE�)�Պ�\\,d��&�(�������b�Q5Қj�VY���<�ALQ���D���J8��LV�}��+�'�ΒN�璡5Q}��
��
�,l��[��klWb�H�h�Qc�Y��l�t=�ղ��//3U!�5�nL���+�Ym�&�z�"K��KG�_���i|�?S�,�*�C-�[����Z����PM� ������)t�a���v�:
�S��R������o���"�SC6� ��W 6�<�i��Wo��
%D1�'�Ӥ~~G�pe񿣃o� �h�� E{��9� �_vOh@0P;����-Mʚ�K��� Ô��[�����|�U;�'�$\z���Y} &\������� �z�}.Z���в{�.�=��1�`�p�m��1�8��B=8���!4<=;�(��)4l�x���*qr��ِ��2T�;n�G������<��ܾ����|�s���V��#L8��4]���w��N���6�5'���m�n�t#��u�N��?E����)�{�v���Ig0����Y���ۃ`�<a�qa� ��!y������k�s*BS���c�����e�D��ȍ��l�9L���	�:���SC��_�Ѡ9���Ɇ�M
��f1�i� �
i�{\����&��bs�����`�vԈ����L�yΔ�.o��{��Kʧ�B��K�ȥ��U�����yM�q��<�f'h!�V�y��*O�-c��f�x��Bvc�|��#�+̳��o�xn����>#��0�GrmgM�
Htn��	W���i�8�\gET�{�@b2�Îq��k�8눝��Ì~�T\>.RA���n�����?!�v��~#�DBFX V{`a�V *���s -����K��Y8��9ʦ���*��g�H�m, � �D��Ԑ���f���B�9���{���<��O���
�l(�A����ə�HW�o����±B�k�/����c��������'*`/\
4!��s0eз
���G���N�*���g�����k�O%d))-6gĎ1S&=WN���Z���@�0�PCP��ƴg�E��&�&�7~�XO�3T�1EθM���~����.�s�=p�0�&����+�	0�N1u���z`������i�^�Npډ�����ư���d~���5�o���*�-�R��8ak��Jy#�ؖdp?K^x5oc��n0Jrz`����)-�j��Z�Ʒ좥݇Pdǰ�X��N))Kcjڊ�c@��?O�J�{����2�ސ-~�]����Vt�f�<�����T�d���
_�?������ն�d��� ���n�أh �(S�7�<��<��r/T�!m���n�~݁�gJ����;jG�{�G L�x����!ȱP��8L�����o����gX/{�%����OL+څr�Y�P���F�!��u�\d��`E(toD9� �t%.�v[ʄj+�������Ռc�+��藍�z���9i
�
�����O����3���7ݽ}��Z����'C�����DB����#Zl&��gE��Şe�ΐP�	��M��_�A�h�<c���Z{��z�����s�I9���gވF���f����N�/��8)HZ��`�mᆁ���-gMd��|�qn��r��Ki�/l�b+��6.�,�SVd&�/�C��e��N�L��U��2��v��MKu]�cӴ�*�������d��o���S��B��S�VWo������P�5���x�]lnBua��~"���Yf xo9e)����{ʘ�l%e�N�[��X��E����}�g�i�_!] ��d��u����m}D5�w�R��[�Z���9/5��t��O�g��S����+����Mtd���~d
tX�9�7(�-�XY,W�"��ND�o�-��}~�'��c�.�|N�SI+f���1���Y�#	
�r�����P����4	]4B)2������5�+Qk������l`�0���0nM��Z+-s�Z������ ���<�����7oN`Ġ\H��1��k�Z$��t7N��l�5�^�ѽ0x�a�X�e(�M�k�s�x
!<Y�.��xs9pK,�����*����,��[�.G���E�4���Έ�c4�����SoP���Ǵ%��F쥜�t�Q�H����1�Vbl)�ڹ~?�<u,�����C7���-��D�����ݔ��"�А���'���i6���v������Q��#�W=��y6Ș��۲�TZ�s�/a�����������u�;���C/����ra�����Q���z����$ڔ��YO6��>����c�����^�$Ӄ�S�����(+E��T<�?
·(|$~��SyRp��B
2�Z���l� �7�U�Q[��C.�ȚE�����"���mЅ|��|���楽��>�K��.U	!��	����8�FVը5A5X�9<ڑ�}FC����Ď�����w�%4>��äk*lۛk�:+~6���LX��� ���ب�$c>��)�?�/�D��l�hW{s��fS@WÖ?R�D�K�eEƋ�K�Έr��[a�,;7��`[�8�>m�Gʆ�ٷO�IQw���6��4���%�+1�����)��9�+`E���`o��j;�V��!]�%}�PN�l@D�?��(O�L=����	6���C�F������"�o�M	r_S$�mb�$v$L(��ڄKN���c�E�Zd4��Tٕe�X�<q?�#��Y�fd���C�?R���c9��i��[���B
R^@�Y?W��k�"���0������E1T횤���֔F�b��� 5����tV!Zʹرv2���f
d�4;�?�_ w���]D�z�<K;�$ �Z8I<���'�c��ޏ������'�Y�����ZJU�۠�Vf���!9䜗v���+�)������7�Y� ����5u��*�yyW���0��p��j^f>���r�QW�8^�����#����yy1��� Q8Q�ň���3W	�׌�x��D�:W��}�^IS[�Ǯ�+U&�Ib����K�߫�џX�fm��X���Rw�"���)1>�u���~�ٜ,�T���q4FIɘ�s��^��	+Ȗe|/��})b��æʟ,3�j�`�Μ�R��K�wU ��-wv7r��ԭ�S�V�d�VOvZ^��THa�/c�#�'գ�e�--�b�d����jQx��P$��NcggT���ǆ_����W=�ք��s~�������2d��E%ԽM
&�~�e���y�����Ϳ�x:6Һ�����}[�W�P�u۵�B$9H#6"o��n�A]�M�M�;�R�����OT���2��Z(��lǱ��^��5��V��>uyO	+Ce+�^]�M�]{�5�pr3@�yV�iq)��A��S��k끰���.�ܣ��Y�ސp�7��He�p�(�Ķ%���ʂ�uɀT������#�:���?�PFс�D,=wG�3�#�l��9�˺�3QlA)mU��Hn	k�#_#kՉBP(dO��h@�S�Ml�y�X��˸)"���ݒk{��7ק�҈c��I��cc�AIȉ�1t��>��t�H�ܘN��̑�xɱ!Ȏ���ظ��u���ow��*\�4�6�\���g�S1����9VMc���z����p�}���,\�k��l�عaP�Cm�>�����a��s�]�H}��#���vO����Q@���H�U��h�&ظ��25���c��2v
�(�W�v�X��4��KVu�BcOU�%J���%�rAL�>��9�G\.YL��`9��Ĺ\�C8�Z�4~�����K�
��eh�W�*gL��݉:i��޵5��A�}���z��6I<%bT��-��>�Q��iI���D��YJA��ge�r ͉�1k��ꕅq�5$�<-�L���L�����&n����K�q���z�����3vhP�����$+�56���������?4���ZVG'W7h,X�cN�LgM[������F���4>�
 (��h�^��)C�B�)&6Č�?�[3Ȍ%��iN.��һ�I-׳B�L`3�_|XeA���m�Σ=�U�с3���D��\<��no��^>�(��x	���T�m_���]�_GJ�c���;44��1��CM���	�Bj����e�R�H2<���	�~M�)|G��~��#��A��正Z�zWc�2j�ݙ l(f�"��C3�ȅ��~:v��j��!L���	sE���l:kp�	]�X����ܞ����S�����T��*�u7�n��4�*!�_8_��X�L�HTw�+}9<�w=�[sUݙ$�ouv�O0E�y��RB��Fa��!Q\�E��y�E-䰜�j�w~���
��{�B�Fm�b��hzp���o��W�q�j.����n����)�%  3�˹[x��N�����'�:輥8��|A�%��h\��r�7�l�>�Ŏ�zr��w�p�j�]�8XC�3�"H��12���B�@��R��Z/�UN�.��x���(L�PJC���H��g{c,�sW�A�Κ�Q�#ݛ%��f����`�'�PjAP�mȤWV�._�,�2N��z���X���\�q9����;Y��R�z{�뜰�E�n�My����fR�ET�g�m���Wfm�Ɩ�B!���48z��w	?��e�}C
d�mB�������vR]i�?K��WN�S�*q�9��_<+�KB4ݹӃTV��TS��j��T��"�wVMa�I�ε&x���ѹ�� 5|�"˒��?�E�m�vp�o\	����䁥_
Ɩ��6ȟ�U�P�����е�{O�Ws��	8�8��{�������JZ��,Bw29�Q��Ѵ|9=c-���Q��1�!�.%��v��6%�=�>�ޣ�Y�s>�����������gw�h��\c d)>a�K��)T���ѪQ����z���E�//���5o�45b��{>�A;Gb���
�v��6��F���\����O@SpO�>Ԛ�$c�cJ9�0��̑����+���/����"��;��K��)yNy�֢�l���3�+��C�����}���
��!�$�Wu����Ў0� P/��c�$S)��s�)��C�MF:Hr�~E:lе�B����i��2!+�5��1k!��B�YWW�	�I>B~�Gl��=4Țy��z痚�N1�^�#-;-tϊ�)����i�>�} �)�_]��p@O�%ׅ/����\��q��]��Fd��o�M��+��׉[�6���KRm��5x�+�����aȒ�gH����h���r��U��
�
�؝[[�!�=1K��u7QP�nFi��^RȐ��C]����mU�w�:�bb��_�f5���i�]?&���Gȭ����j�ūq-d(�Q�	`�p�K�A܊5%D�\�P.�D�>��ZADYN�
�לց^��;�0-;&h�
e�L_�DsKר����=�Z,����4�GO��-.��|�����@�V\�>2J�t\>F��4���1�4$��k|tm�j$��OL��I*�ƚzS��W�#8P��m��LG�&�tU�	�[�-�H'��V�4�j=�²J�O�&��X-�ƴ
2�<�3��k��O
����Pa'�"Ƹ���W�z���l�mi:��䵆zz��a6D"��������v@���j�<�KqwV���y�ɔ^,��S�rY���ˢS�5��6�9 4���� T��mꉥ����1¶O2��Ę�ϑC1N�Ǎ��hx�����+XCQq�1����w|qE!>�%�A����t;/Bpe[y��ҕ{]w&.�y%�-��W�U�xϺ��Mv�c��د��⿇�n�ܮ:����.ݹj����'��2�7%�Ŝ ��.����_�J�,^�(�������#.iX>u]��8'	��)�fE +�.�/�~�o�c�!��_��0bp���bPSX�=e�7jæ��j��A�n'�lm�����c�s�feN�yH#��+:$�����2[\� o�l<^�0,e�2}Z���<�}6��%x�7�^8�ˉ�� /��{�R\bZ�|�I�ʫF?2�����ޞ��wc��[��> {&�KD�̱
�"�E�:Lfz�ty��f6ɇ���pE�[)o�,	_m��MU�/4����P��&
�L��N��e���q:�g��p�%>q�
�j�����q�%M�~��䘍�����l9a2�I	��W ��\d������=�����8�\��',&͏��.����U%�n����{���ӗ��eT~�=�E��_�{l˻�^��e�*�
Bb���H �sYis�ո�� �<�e��U}/U6E�"���n�9>�>uC��s[iXCwZB��7X[^�AX�`Q�xf�p���&�U�VNfʑ۲g�\(9���O����]�9��~_jp���Ͷ��[���
Q�(S��a	`��ç�X��S�М(�p܉2�m�b�3�� ����Ӌ1K6U��,��.Pb�rg������5�G������`��A����Okq[G����am#C)���,Ĕ6�G >�cn+����|r��m9���ǐ���&J|:�HV��1�!{��)/q��RQ�=N's�ٹ�ʓ����������k���5�oG�H���Ejz�~7_k6N���(�S�M���_�'���v�޺��I�e"��_�n)6�������]��ས(�5����y��VW�"����Y�ߊvf7�h�T���֛�8��5j�JV��7o���$��Sގ���3��b�ʲAv7=�A��Q#6�`1.��9p,��=�}���8��j����OC��/�D�k���q��^�y�x/�֑Ev�)Z>�f�I{/���\�qm�N�F��*~.N�QT�����X�S�gT��ȃE~ë~	����K{(�wZ~�\Ǘ� dP_n�G��� %�K=Te�����
j��V�8 ԁ�4�l���'Y�e�#p^:/]sl64�؛�|�_Y{�ht�
n׃�&J��+��24�`ˀ[eD�+�#BZ/3�A�A�y��P����fa����D*��/`-1k�>�k:=��>�&��Y>$y�O�{��Bl��z�'���o�����侴����g�Nl�*ڥ�"_�jؓ�"ҽM��.���4M��w��l@aMܿ��'$h1a���!�c]HbNz1�����f�@����{��<.D�JU	�*�*���w�VD�S27�^I�%tE&�>i��:�h�f4�{t�)�c]�I_�Ѧ��+���wzG���������$�oNWU>[[���xt�@��Ŋ�6�+B\2^��Uy?h�y|F�M�+Mޣ���$v�������u!	���Ys�~%�MN���TK."���Xf��#m	����yRT6i����&ʍ��Y�����Aeu�����0���\�Nα�������q�XI uY̫(8u�*�us�p{�i4a�h�jci�V�I}\��CEcx����'ƭ08���}F��ǉ=�񡓯����Cw�8��=����+SJ�Ǜ�f&`f� �v������	��ą��
�&����6����0�`�L�2~d;���]�3`�N�]O�Ǟ�@>�88�c��C'�;�M����y� ��&�����3�Pv̓�'O<_��<�Fw�T�lHW�j0�18]f�����T�K��-��5ŕRb�2�z.�X�	V���M�)3'4��Y�y����ڋ��,����j+d�[�L4M��8.���\�-�C�|��D��;�ՐN��� ���V��k#Jú8�~In������~l+���x�Wˊ�t�s�X����a�^w�{LO,��b�j�۵^d\��N_j���)��`PP������:�^���2gY^~%��7�{�~v��K��~f���a�-'p��g�t��2_HX�Q�-�<��/��Ș*pa�n��5����I�`{�2)>͓_X��:���֜����+7w��M����->y�a�i�R�^_�-�F��b/+�|a��|�q�+���p|-�
���Ҷ�i㝫P��PT��S�;j@�(T[3��\��Ȇd��-�1^����{�������b��J~>x-8pd�^�Q/�PNy�W����ۈ��z�wbE��56.�{2����3@zubh��J�Q����}�؍81k���s���Ief`�e /��!O���y�e�9|��O���st��|&�a�kY���ݔ��uX���4�!7,#ޡ��Y�iJ(�Ϻ��J\��g�!�~Q�U���Mќ1؋��<�D�N��o�b ��a؎* ��}�Ƅg�����|�4�� �Q��K�7	�ZR�T�p	cj�b��Ik!.42�?���%�0� l+���/x��:���V���(�IO�Y]u���o�%	��f�('׵�M	 7EI���a�����Ybh����<�oG��X�7ϔ����o���ޭ	�Ըu.�D���L���A�\l0o�I���Aj����0���#��@=����P�&�Y���sҠ"5a�;��X8/yE���T��m+]���D��*�j��$�\��c�qdQ!�ε��rku'�`�9n���*.d@+F���=~Gq�Ͷ�����yEh�#I�8�0=p�V���~ �@8<�%�Mx�-�;����$���`[T餟��<N�騱���-����>����XB��G�v�����(Kv��sJ{QcZ���V#VS�ll�S����i���*?	���=��0lE�}D�S�4GJ�7~��4鳯�N��5Sʭ�)w��*��ßɧV�삆D���~�(�� s7��dո�Ц�� ���!���+�����@�r>�J�c&�gH��ɵa��8�"�y.��9㙅��^�� P���?{�k^{Y(����$�|� �G���i0!�F!�~������{ed��Eօo�t]�~_0I�uǣ�P(k]S�gJ�<�'c� Y[Ҳ���k'�n���1�38�h���@���0�����ݬ�㣵Ԟ���=iKB������QE|8:��(���s�`"��7��:0��9i�W��CV� �m����?�l7ރ�r��\,z��㻀��e��#�Zo���>��
�oI��>6���E��B�*�fOf�)ZE�v��r^h���5�^R�vQ�5Y.'�ɰ���ڐ%Z:�l9O�	 �Q)C�4T�_~���\��Al���"�������6�ͽ2_���?���2ӄ���^�bҫ�	��=��8�\3�[7Y����6O�g����F.D��Vx�:ܱHz��Ĭ�^|*���@9�AK�]��&	�mѷTY�`W\��O��~Ҽ�����0C�s�>��4�x�5�K͹!od�*:+�CR�L ��Gl�*J�ɋ��.�=��Hup8�}�e���S�+W�dk� C��s���q�Lr{w�%�k�eR�����O��ZsK\�r࿴��7��Nఙ&:76q��fH9!��s�v�G]?t2�8P!Q3��΅�clS����($%���D'��E
%bW���@U�Z�F��#������~3��vJ9��RH�w˖H��/�������ß�*��D�Ӡ�p�� �L ��2����ri���{dj˒����@>L��$��� ��\�`=�L������&DϺ8{@���		�Pn
�t�R��N���/ko#@�ć-ԛ�� �7�JKc�B��a�:I;����ʮ�4"h�K?.��`�ۥ��X��Q�&ffC&�r�I*�V�f�=/�$
�:��,��j�������^���J�/Z��Y䝝�Du�w��� h!�h���х��)�����/&'w�6��W�˯D[��fip���5�]�T�Vhї�Y%Ҋ�Όi�¼j�����+�R���t��#P�h47�J�L)���C���ݽ�A�l̻
O��_�G�"Y���w2W���)�H�{~r���<���}PDB��� ����`C 1��MfИ��o���K���3�@<C3�'�h���UF�3��x\�!�z=1m
�#}��x���j	Z����;:ğ:y{%t�e�X~�ء'�aI�
"�)��y]�������z��<��5�6�c����@��R���F�?XޏY���ˇZ�f��`���j���1�>�_�V�o=zD�֯k}�Pm(�4ZNN1<�O�&�E�� ���8tfR*��d$2���bc�h���R����ȡh|�3̞����/�&��?v��`!E��vunzb�[�v���4Y�Ob��>xܪ[Q|.GH%w:��@|ܗBU-�7���Y�ǫF���R��8�}��9z����alΟ�{��Ǹn|8󍖀yP�3jJ�ݑ1�"��m�pO��^�!?�6_1Y�I wyzgP����oS`<Ԙ�fA�D��?�eĮk����т:(���)�V�ˋ
H�X����	
�U�5JJ/���¾�9e��*��;���猅�߁��7^�(6[î�|��1�?N�xg���߫�z��	0��퐜 ����:�[�o[`��3_1�7�*q��$���i�:���<K]ma�ۈ>	�D5��PG_��v7o�>�^fR�����J�t��7����@��� ���/.�O�fƭn�r�Sɨp�(��X��_�&�_�������.�<`5��,~̨p�َ���y�X�A�5M3c(�n���V��#�HK����(�J� �ϸh���ş㑨��C@��{�>�%���mBi�r�;h,�T��Iͧ~�qv�D�8X\f@&�(���Zf���⤃�S-$%�"��b"�[U���^F���X�Id�L��tO~S���*|�#�7�sD7[nx#̺�?���D@f5��ƈ�F�ܴԄ�X���ݲ��(o[)J���$�^Bmc�������K��C������-�` ��fKz��o��1C��)�̖K"���%H�Ѽ�K��Vu��%�@B���9�&���H�+m��;b CٴAq�H��j{T��oy߂e.2��YI�u���#�\F�	�%1���4e�fHmy9Y�F�T3Q�07��4/&�h�tts�K����5���3zYr���2eu^C�~�C2R�2��t�/�7����l�S���}6$�E{�±�����c�X��Vm:�f�E1�Z�j(F����]5�f��: Xpך�|;R=&[J�MuE���$��ŷ��J�!9͵������kK�Є���DY��Y�!���"��dy]��|���{W�����k0�О�C�+b1%�Q��3�vaG����)}�%����U!#�V>f���q�bsK��!��`]�4t}�K7q��"�ěܷn6,���=�C��Qݎ�G=<�n�sA>А��6t�"X_(�bHA�����$�..���E41�����&�������S�A�ĥq2ϖ��i֡����$[����f\�W�ww&���G��匒�Ք��bX3&�5���%ut��#u���Z�n��.4�x]��^�N5,Hl|��B$xH�B��������n�C�U�Ȳ�e_��TXD��R�C���I
2���ޣ�pB-`�J�/�����?�]��l�����)�٥�X� �f��z�s��j��3鄔A�s�i5XA��1e&d�+����VJ�Z��Ex���ůc�71z��7D�j�f>^���Z^ .�0��V
�$�l�ct�2�� �C���5"���r�١� �2-�#���#��X�n�UYܥ��:���3o5E1@?���{Cje{�6������pBf`�)��W����&�Ғg��e��I�>^/�h3�}̬�v��,�
p�b6([�1bri3�nOsѣ_ό%J��U���p��v+6��zs�gi���p�s��b��Oi?�w)V�J�J�S�э��E��~i��V-�"�)kZ��cH��"�	f�釜�s�a��;`
t�����]�[�.I�9Jw�X/8[�q�RVf���\y�`�5d����W��@;�m^�t��p+xUݕ�z0R@6;�>�G�t�J��,�j��<ݏ��q��ܽ�΀�,G��OH󐐾���`R�e)[���?�O�w��-&Е�b���4���m4��s������EeV����s*��f�mo�3'��wXr�A��{!�\�Q��H;4ߐz���MFó��dw������"ԋ?U�G"Ħ����*9P���O8�B�"���Ղ��?;��$��W�i,��k����	M�Q�`���$�R�i�d�L��<� ���w��e~�-C.&t�;c��&�8�~d��o͌�hΫ�:Ν�d���x�C���#�u_V۴� 6����*�k��Aq{��% 0�wA[w�)`Y���8Zn�Ђ���Sy ]��'%=�FW�)S=����6e�v��_�\mfE)��J��1����
�'\��vM 	6����������%�ާI�D+K6���Tz	����n���-�Ȃ,�|L��r����i�,��ݚ��]~2�	[Di��Li�2���k�*1��Murȯ���J��4� �
�;.��C�rĀ���r9���|W?>
��C9�yD�N�T
�ͨH������bp<C�a[Db���^�����g�T�.H��ʘ�B��v�e͝ŲT<Z%��6���� ��[&���P����O,^���!z"=n��Q�G�y=�i���_�ySK^w�Y�a=bm(����4{&����x\��	C>B�Mx���/����q��Q?�t
<�0��w�;W�cZ,"r��gМ�e@%��p�:ũ{��H�:��'w>���N��a�@�|����Ʒ��ш���n�ͅ9j�n�d��G��8�U`1��F���kq��<�c8� *H���&=�/��'��eW���r�R w��<���5�&�0e��9���,���,C��a?�!�ϡ���R��B�ˇ�"�����{rw��_M���j��H�ӆ*�S`����dq��_7��� �;&�KxC:5�!��btE.A/�,;{���+#���\���,��)�q.��r}W�b۝�1���n��Cx¼}��(Nnxo����y0nf0<�w�U|�J����J�D%&.B|$����0y��6?��z�e�v����pW���q��S>��^T@�9@�Ι$o��j�(|v����z�>Nc3�F�r��B*�w���r������h/�|G�����>5(����^�7.��!M����q9��r�g
�i&�"Gg̰�(�����)!��`��D�?&b����&֢Ӣ��^=���G�z.%mu�X4�Y���5�-%�ҹ�IZ���(	h�d�a��P'�U���D �KֵH��O��+s�+ ����wX�)�	�垀�TU�O�	��m�Ш�7ے�g���衒��v��QO�>{�/�]��2��gf3i���|j\%cI���=:����y���d��ք�"���gf�RB?��Pn����[L��H?VƩ��."*�ݚ�d�c��(�C��a��}T{�K`u���}�3$޸A�Б�p۽�S�Wǿ��W��������Dq��C��__X����C:�$���������u�}jmt����_2�����AK���w"�yC�>�]V�����j��-���a	k�<W}�f�{���k��1AK	�H�R:?"ФE|&�e�>�`�yIjAW�NQ���X?�E�4�_�%��bD�l�^�Ej��޲5Q%�Q!��Ѕ!�#���ȯ��� T�*_�K��U�WGxjO�-E(����r�o��x� o/�'���S~���K�%[i�O�:��e�Y=b��H'+	�:IJ�ɼLR1NTi�Ǜse�n�BXБ�U蒭�^���(7(��t�X�jiBfTO�l:;��$ehC���B�pXl�H���!��j��4�#/&2�ĔOD_�n<,����O~R����z���(��j�N���B�=�]��Ѩ�W�{sW�T`M�k�A�{#=��hF�h���X<�aj`�Δ���|@�G;�bP��U6��C0���6[ຟ����� ����3�R�WO�o��-e��jw)�x4�m�F䆖n��
���`�zA��R��`lq�OS/d8�1��7)rs(md|������J���6N�&�Kb"��A-��4T`�n�8,�F֛J2�[�NG����';$��
 C������6N,2!�;}*�]��AD�ae6�;eKؐ^�����U]gw�I��
�_���_\�=>0I��!���tKͣ�Tf��[��.�>9��3��,��/8�c�F�;�oş�$�Yȴ�M]���v	�H�L6��E6q:,���F�a^$-/��Hշ�Z���ӜA;��@O��~D�n��8�aK���|k��Ŷ�La̾�w��+(m��ҍ�df)�����Ž��X���Q0�-2��y#����V�Κu�ښ8
Yॱ*��΍3�f�Xn�[��o`�N���L:TS����ڧX�<BQ��]v��� �"��NVx���[��Z���e_��]\�9��n�3��/*�(u7��~����0��s��?G�g�rnk4V���=ݿ���z	������}z����v8m�G{����;7�pr:AC���/Ә��vlA,Z�+�����ftŠ�H�45
���^mp�ѓYd���\<�Q�Uy�3�#~�3���.Â�t�eL�L�v�F��fb�X>!P���eh���ϷH�'�~��=�PD�"!:����u�.�#�U'	�]��Y�ى���''��IS��f:Ƒ��Ԯ�Z]x�|�*��FZ�w��]�1���Xd�L�.��n�A� ��(��R�������]P�\���lE�zEm��Q�7�� M���Z��A5Q5�CFtuv�G���$�Ă�|��MN�l,i[��#��Ub�/rv�S���dW��U��~c'��O����O��vn�V�q���2��;a��9ݭ(�W
4	:⾽�o(I�.��g'~�5z0Mp6����0t�w�Wdt�)�cV[>�j�"j�������W��O���pP�I3���Q	`ը��"IVH�%����2S��zJ��������<Ҿ�g�И�0G��I��J����n����	��U+l'l1��R�N�Φ�����C��b��>�~�WKd��DO��\)E���R�c���u��F=��7���ڗ�f��I<�+f]	e���N;�?A��k�D=�[7�����=\4	joi�:�D�A���nf�]� ��d�u��xI��v�]:�݋���KQ~�P7�]8��~�l�GhH�B����84"㥵9L)|S�I������v��A��Y�&gt�h�����N�P��/�<�F�O���T�,����1�A��'ػ��C9�E�N�b�78|&�k��pd�e�dt�?�(Y�a�H$1����Vu����RY�,ȝ6&r����v̬8������5��b����k�8!يc_�*�v$�&1�v���&�^���{���&��(�p&Z`��Ma:(�	���z�W�wJ ɒ���k�B��� ���5�Ly�<T	�d��M�K��rVoבn'����R8&sR��ط���P���|/u�q��s�u�Wj���ܕ��	=%n�N�g&w���΃k�آ*���5;��d
������7�Ƽˊ��p�ܑ�9�g)�>x�.kᒳ*�Ӵ��%0!�*�c��V83
�5[ :R�����A�:���+��;���60[��Mr�1��44���A-���=75���r��`]�5J���_g�C���)�n��ӿJ;rf��g���.�|.Κ>ϡ��P��/iV��~>�\����2lK��<��$�NIa���/�ڳ�3 ,�7��T����3�	��o �S������p�U����j(�"��]�_��׮!ټDKī�V�s�P	�aP���v:^���v��@/��H������sڭ+����EQ'D��ضb��H�|�x�������?���I��������W��E�Z(P��#�=�z���.�X�l*�l����R��SN;%�C�� ���J'[z%3u_�D=(��Kh�]�|L^0�N�i�i���.B�th+�a����<zssv�N��?��岠��rN�S.8��V>:EyZMW�#| �˖�+�( �7��N��O�i��am}��o�*��);���B�V���k0?�/�8�{*����:K�N[�Hh��i�zĚ�7�ٛ�P��G$�:UL�>Em�Qgɇ`S[<r���B"mž�m�ѫ,�H�Z$���wEr%�}J%y����];T̔�=�����K6-��� (�c{ �Ϩ�D�����8ȫ-D@��~�M�Y �~��B�U����T_�>θݨ�/"�@�]�;S��C��\���
���>�R�·�&7�[�[B��xMho��3�6�u���R��	�)q�L�����9_Lq�/Zߜ'<�9��5��f�Ũ�͢����`���&��\�Q��+؅��\�H�*�A9�����g�@j���L�mR3I#��>_�dG��q��s��=�V��t��� {���!C��v��m�{�<h��&:�0`γ�󃈬�]�t`�ǃ�A�ؖ��hǝ�]�r:��k�0O`��<�NWD������x+����ץ�����9�R��`��aA�z#w����#��@6Pj
W	��>ޜ�G�A�~hZ 9Kb�y ^4x=�?0���Q������7��Dd��o�QeVT9��;Y�Sz���hA��Cs�[��Km�;��EzXJ'����ϩ�8+���+;�Q| J6�L���H��`c�L����ƙ�|�.�l����OѼlS3\��S�l�dK=l$\�3�ؘ�0$��S�ϵvC\1��u����ݔ���U�(���iujF��Kj�U���т=ރ���|A�����Q���8ďUN�k� 'Xz��E�4y	�F�#B6`�nP�ߣ��ٳ��JtĴn�?"�l��9uV�D9w|�x��;n�h����E(�?Z���������s���+�kV��"�Y0)���ȴXj�a�O{j	ِ����*~Mǫ�$��������1s���V\;6��YIߨְ9�vo3#�
h:��]�R���ܓd���݇7�JO]ć��� �	����k<4��9��6�т5�j�v��b"��֔���	���A�&�ر�9���v)��/S8��0�"�"�q�5�"f˩�9L�k�bA*��I�;��~a���b<�cn�	�Oy�>�5��!!����/�|��Ƒ5ʟ.��)�}�����/)�oBmd�6��]�i6�7P�@�8A�
ۚ����{"��[��ؖ P����qՕ=�bR"ɓ3����ۦ�J����?	�]GK��B\)�<0�FCy\�M=9�ҝe=y<���"�~��V��y"�!�P�>c)�d��p`�R}оP��U��|��8�	��Y��x�	�;�V��!ah���D��>��c�Ď������%�zz w������^r�W��\���Y��n���S��MN�ES�s0���`���z G�& �I��#�9��m�J�4������Y�M'�	~�	��}�I��m�\Uu.���8�
.���iV��.x# R����s��I��3��}xs"�B�LG�HW��.(ɿ�����*���V�pW�Z���}�B�g�&[!a{+5cj��\�dCy:�%�C��Nl.�����up��m�`W�z�yAi� �_(�NLQv�|"��qGӂ_�%�؋E��9�f���엓�	�@� 4�)o��F�G�!��,fN��Z�>'s�:�N���3�6�[c5�������s��g�G�����A�j�E�S; /�}���A��U���I��,�t��u�<���]M��-Ej���D}�lR7�̄L�+JZQ���9ro�[g�ܺC����(�fk����|7{����~p�����a7U�&uoa0���Ufu'_eVh�>$~��6|����9��y�T2'A�-��P��rJ{ٰΫ\%����r�EW�x)3Vs@i��v��RKR� {纐'��?�7>�[j��v�A�j{�ѓ����X��dnz�sv��!-<_u�tj��2 [�,_*�S�n��G��'̱�RpN�nݚ&lw_�{Ӯ�ZgD�����5��l�%.]��i�2��fe�s�f�nc��go�X��?� *����E0
 �>N�z�oS�`�UГ��Q�c�zҙn\68��#�.�Md�!܏$�\C]��:��jPc<x��d�9뱓��>�f���~|�4�j������p�2D/��J���!����z�F��]3�E�l��+�SH՜J�C�-k�?u n�H�F���0������|c~/x8O�N��i��T��
K����>��a0j�9+�#,��+g4G�YF�CW�Fug�x�LPn??f��K�`��hܡ�ח�GwyJ2�,�2t�[�.�luq�|�!����mpj�=?��;*D��)\��]��/�%/S�5yjqk��j�"�u�Zz�%*�b_��� ��Y�^�	~���t��-�؎���B$����b�aDf��F����m�	����x;��(}�rc]�{����2 !�T��z��N�E��>�y�y�EX��k)���T�ei˳��7A.��Sz �%�
PzX���k"7�" %����T�Z�B��=t�t���6�0CC�����7�g�������!p���,���*C�Y���̉q#���VLLg����0~�U�ңO�sL�m��/$}�S�,���ftﻻ�j@�O�b�����aYpK�r�E������ÿ�Ћ���#,т�E����E����<;1`�6�+s��X ����G0�G� �\{�x(���a����	�jK�^݅d�"���^��@�b�N۷�x��q�����.��m7�`@��I?Q �6��'+��t�b��l��w�Jo�?Xa����u���Q�^��q��ƚb�7?�(A�d����H���I�0�Z����S"m�	�=��-��F���,���x�
J�#�2�ĭbFM:ծ�縁��z9��R�8�l��'�������MgP��{�u�oe}�0qX����zB eJĒb�en�Mlq�#R?�e)z?u=��;ć���GLL�?u��sA�[���>����:GA�˼��{�Һ�k��u����1@o�^!yߗ�bz�-���UI"TE��u�X��`Ǽ�^�vԌr�=I}U�B���A�ф�?Y(�:,y#�EY�OE�}��5	Q��Sff4,�1��U�`���tK�`k�	�Fp�NYp�Q�Z׋��<3��P�'����K���Q\\#������JH�Y;�$��D�y��y�?��u�a�,s���i�O�lؗ���&�jy:��S.�4(�o�]ˆ�
:��e8 ���s���si�����O��9��YXo�7�}$1�{}X�6N�s�<�a�U��Sw}�,�g�Z�:8.PH@V��ԧO[��>ZF ��t?�%���h�"$�	o�9@w7a��^�eSH6��^o>w��}-�6-6������c�e��8	+����Oc�駊�7U��� �D��1����=̛��(L*xX�)��Qs� x� �#��\`��N)�é0�$$��S��aB@W��qA�f�W5pF-J�����L�/�],A�/{�Q������v���'� �By�D�`u�*�!k� 	�`B�㝫Hj��E������8-p��%�(3R��{�w�-���t;�@�]�������d�vݪF�Rx�@���l3��#�1O	�q�Vt1�ۭk����wN�c�ؒK1-v�`ͨ�YaE��h#׹y-�"5@���J��8�ؼ,���#P+ch�g�-,�N�o?����Y�]L-����2@����fcaCU5�U�r1;�A�BHS\e	�qz�h�fj�L�~
�B}z�x.
p��q��I)Ь������}A3�G�8ۉ�����l��0�t�ʸ�o�Q��71O+�����F�L"U~+̄~����ꨇ@���'P�U���5XSo�VP3�ᗴ���.X4_/�u�c��zC$���g���/5��hA�a6D%�a��v���4�{���a��(d��jV������ުT�]�P ���j�?b�&�r���D�(���a�LhzHK�|�����t����iM=ֿ���U!��6ތ�hW��-��G*��9Yz�H0���8Z�-D�Y!�s��b�S�IM{I�A�����0�[7��^D���A !s�Y�PN;����5a����g`����JGm}�l�����M2��q\��cX)PP��n�!Rڨo1)��ПSn l�:��hp���[���3�N�i����?�-�ҷ�ǒ�����}�*@��OC1
�ݣ��k�J����\��s��Rǲ����*�SA��a�U!	t9��w챢��r�wbcny��H$)�cQA���D��eF!�	S۝��Z��ȅMj,%�n�n�[�6��������ր�j#=����>�iS� ������Z�R�o�Q�1��'id���R�ځ�T�Pq�%��<����@jg��l����N[���Ҏ�$��)_gcF��C�O.�_�ŃO�fl�p�'MQ�u����^�G�#D��;�f�3gs��k�o�^�!���|f�A��LƜ�ORɍ��e��G?�4w�I4��D�b`�����b2$�4v���,�EO��?}��F�.:�����H����A�4�u�p��
��k�!��!�'����GW���6}�pl3	o��Y�>V\���j����S��C���s�?fF�/�f�]ҭ�ǩ�|m/ı���ۼQ� @���D�E��&�Q���O�ûn�i��3ܵ�:��_�P�9ɗ]��I�Q1WL4�K'�@���c�)y��Eeï5r���M����m9��g�A�ڼ�K��͈�����X�lD"x9SA8���� �w��f��ph���gY0����Qӯũ�n�
�fMDBl�r]�����Q�2W���bv��G�~i�W����ȌR� ��4��jm�?ގd=����d p;���t��J)餼�V��͵�H���:���HVN���̠�������q���t���L<�p��'����B�}��!a��f(
 ��1ގmu��`%�ܗ��A�H�VH��Ѥ�[C-�:�cn�z=Ti	���/��s���d<�L��c���wB�h��J��:w�W��&�*���
�,�Љ��S@�+E��(�.*��4���$�+�q;�\�[�'|-�������_i��a	N�ZBFqmA���ȄՎL�^��[O�~���";��B!˓�b�;Ck�+�UB�y��W��[��$vȑ~~�w147M��[a�Y�O�_9�޿�da?W�Lr��k�7?,�>�U��QQ�h�p��-ĳ�̛t̄���H�	"��D��^�����%�e+�`���7���"]�eM��,�5�M@0w�䒖�&�"�����|gyB�7�[��j)	׉�S�'-�Mr�ʽ��Sq1	\ٴ]�[3�QJ���Oԙ���1Qd���k9�?a�<y�?\B�q��
��҉�}���e�OK%��a���o6�[+�{?ז:�H���0�N�Ij4���߀i��?��x�����F����i���a0-C��,9:�8(á�a�����Z�z��A|mյ#�Î�g:3
�׵�y�yLșz��`��Y�~�S0��@��Hr�f+ce��y�D����T���i��δ��o�����Y,PqT��� ��5ݵn����ɗS�,�PH	�m�勩z�R�t�Ƞ�q�~�5�sѾ�r��l��l�L�毼'����JW�	����0GN4�0S2�CԳ �����;�2	F���g�]w̛�@�܉BI.��K\�DQ�F9�|&EPG�Y9$��G�s��ޞ�j29���#��f�
]@��몌���w�Lv�3�db���51m6�p_�ū�wl��w.<�c��ը#��[@:������S]5%v-N��d�*u�_g�>! �䞰9`�1�{��=��e�o�m�:���J� J���k�로�p�|��|0���ѓ�j��i��YM�.�cp�;ft��i���$�����D����Cb�0z �2�w�������]��
�|�����@{��@��-�M[iE��˞D2�r�2J�T�k_�/��9���qz���G�@�7dv~u��G�B����RׁtN�w"n�v/j��&�L�a��Z{��P��JkV�X���Q&�s�5Č�"2
�~�_�>k����z}�~���Z��LU[<��!�%%����5c�G�����j�_SªʱW�+H=��R��/�f�L�g&���ǳ}��S�����RtR|S���H�%6p�;9��4�-��|ЉL�Ip<y��)Nd>>�Rx@)âwY��"~�Ȳ� �Q�[�xwd� .=/��rR7��5���{�,=�C�m،�&ھ�%\��0L���\�dܭ�{�5�t�xppB2���$R��������l����]�1';Ѝ9���66y
}EkT<]�{d���n<��?� ����������VU��Z��mt�c�;��8��	#g5ȶLU0�O�����X��'��=ĵLW_zw��.�z����_D�;�K�_���L�"���m>z�O�YX�K��
�����O�X'KI�8>v�ƹ&�Y5�S���^�쾏vO��Z��f��՜�~~{:m�W~+�W��A�^&�Q|N~qL����Y#W�U�'b�����E3���9b;�w�A�t�ѣ�ucJZ��������NYlh�K.}����i;o	��g��;�D"C�%^6��J�XE_G�){�9a7�b���Z�Q��o��n�Z9p|w`�+�\$� �&1�T�GV1$���/�M��~�W��Ð��Xn�@��� ɗI��D +ж���r��УB�OO��Ql��W�]%���B(�d��=�")Ȃ��x�/$A.G��~���d�a�=��r�F�>{u��	�c���5��r`l�j�F�Z苄����<�)���t�� L[���L.,�"�^-DO�v���왺� >�gj�ll+�c�^FcK-�O\e���o
���)����&`�?�e�N�L��L=�t�r ipv�m�ۊX��i�M�HhHL��o�#�[�ЫYY{��=X�P��	�Z�<U]�6�s�n:^N���TDԡo>�$��*S�\k�9@K�c(��=b�su~���i#`�#����	;N�+�i�a(U�v!_؀!��Q�
�ť���@�Q��A�B�q	Ü�e�)�2p�=�Y}r�I m���&n��	���a0������-*t�?Ue�A������
�}ߞ5��k5�7[����+�b$Y.@K��J,���}��p�SiP�iT��*���TY������ʄ��'����h���������ab�I7�?�\�g7vB�\M�)�|n�!�?&��M��]������!59�cB��+��Nu	F=]����Cϛ�^����;3�p-��F\}�� �4�X����F����[���aH8)Lz�u�Y^i��cKL*v)�Y�%�?��a�K:��_��B�I/�<�)�+����������g,�P�;�� Kt��v�ׁ�q
Cg�b��@Y���=ߍQt����|�KR�F=�;G�7)s��c���{*���$�����s�;A�����B����n�&D!�����9�`6r�($��3ܩ������s��;�(9s�O{#`L'=��c1���c�MƔ���}���0��9���w��to�9P��z��0<��>Hс�N��o��"k�A���C���_"��5E$8B�PMX���u�'G��^�lT ���C��2{��N�_��3�z^]*¡�TYX
���Si$=+崈i�eK?s������0�-K�8�CAV%d�gs�E��ylx;��L���������W��  �+kK*