-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
km1fJDDbCF0uPwdwnk4EQmtjp8GhnLdKDgwWhcyl5tixSI9lmcD0qNiDattaZg4GL3XShgC0gyQs
XLPeuN9jr3y5Xpd1iBY3g1E38KtmBhijck94p8Jpn75zNwVldkmUiknGNRWQPJsaF/r2sVkabx2t
LBiVgUiSlC7nLONJyR8RV0Qg2DMxKxlvLfE8z7HSde4tTpkcQsWcoMXbgzEl1T+PFgd9cfr/jQnc
vul03tUWNrZObXogYIWP75ppfY/6WgeO8wGjEQJ0bDIpdJC9UEEG9BVqbA84zATGnqcMfYCOn4W/
3KUaMzv9MVIpulFv1tAhY8IkvCq8psIcPA2ZNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
JjHXKK0c2t8tmsTdyQ4/sdnHA0S8ajox5beFc/H1sOzYzLxcqTg/879fQU1IaaHYN5dPuS1vZif2
xN8YYiyeQkbF4tNEukZm5H32hKbGTqeLjFaF/FCx1SS7HbsQ9tdvzldK5xcIOg42kx7ruBqnTmRI
V3i6QHUDWpwJi6pv6YgAPFZiA0kAXiwnNCfRnQ/Vh2+yYzEyaqL0WZfjVEpQjXDeAfBjl3gl4oYR
tHB5vAgubNo631cpEbWjOgWsNz14xmf+8UUp4JhsquvwvywB7uAfdeVqh6ZBwrPEUBbYR38wOOP0
nrzXUUehZbJKwK08kXHvXWDb3T0+qMzpmd7JlIQGqolMRqtX7qGkz0sPElCXzW06NRH0LhNbCIYC
g0njNHsIFaV5qZZM9KoCw6/CjAfgTbj8LhjKESEbYhZiqIZuFOBmbqe76IroiZhmQ212AAdNPD5S
RVBRg+xCsyIrn3RoyBNIJDT6sAVEXGfqzhPc687baQOVSpmooY67FBYkA4nQB6n8Z2UI7FdXqC64
SWphZTjbvovzt3/uIR0jExGzHfyfK62irA1X3L5BX7D7FlZcd8CakUDHyaeyEat6gok5wXau7r0u
kzwllNTl1j2H7FL4SWtF3jshh8CbiMKAE9hy6cMheInMgpGhka7czMSgz+SN9OQ9BbL/oyLNwQYn
EOU5Yh8oy9R8n294pPffhPttLSQHbzpuXt8K+bx2M442jBLft/lhe/281esZWg2+2QUD/rsDsNVA
/XbnYiaVLq0yRrppQGtWJngf1LMLycHE2qUxzVUk4NMfaYutik5npZAw+SNWpoL4gTrsSGfAnOPC
p0JTHUk4q9LKed55QzBc6fe5GpjFKaM0RDZmzFEvV7+D6qlVXWk7xkOY+tqjmSyYmElMoDuvDIBd
AKhJXBNX3uCfovylUMuDM+1gebaHmBr7tCFERRj8cbEeLSjmf+2mtc7rr5TJXEbhvQMkLYbXljMK
FCET9MIA84L7etzbw5Om4BUByGIBCuhjdsf34FJblyBXE8FQmkkuVhgPr1j9pMfT5M0gdgZifLt7
Urs51nOX7hMspUArZldx1APbjeWbaMaYmbeWxE2CwwPpTqYMrAeIER5/rU3uOIpNEjbecxZYMqQC
OL8AiVdjRurTuJoW1STV+9ImymTzkN6jCehOKcbrEU5Dsw0XQfgy1g1MfMAdQ8Dq+2+fOZPZsOYV
Wfbqgo6ZOiFsEfoli+LBjWbZB44kD8qfNAwNh6hlrOAVdS+FtFbgNkQGL3qgronRCmSM5fxTfm2H
UVe+V++PiKTsnaiMxgl9zfWQJnOtqAJrpJjDcOIaDWEfe+ULlCjBHUCLKP/jFwj/3XMBH3KGgKK9
YUtRjmSmm9GrQwIei3O544RVxmbrCS8bg7L2BLtT0/MOjNIAYz13rdl4bjOSGcvxxUHxroYRi7G9
o6dqNk3wjPjXltSQAqnu1GTLDO0XnVpviYrtUzexUJAKwu2zY6veFGES6BXanif/zNwWWA3hZxp9
ZVRV58GNliRU/IRtNR1elicU3CrqsCIaZKcG2lJgO+X6yZSffoFWDPmC32AAT5y2OEoCW/I5tPAM
ngAgqfBSGy1n9lMlRdDMPUXMOOr8ExKq6z5hVvIC/9NLctMOfnfva+s0MvLKzbs3YK2afIJPpqff
r3jtdmraBUfPxgUNdIc68Y6tOVmJZ6XpLOTOWWwZUv5U4lopdVXfMmrEwtkefIgswx8Zf6KcdrMz
3k9udJ7m7LJKbFelzjuLtMBZWqqGakDaTFv4jJKvsj+bpGN49o5Zl3xRbq8hrtzSLMMIsMXIaLL8
kJUKO3GzINIwzUUjVhxdBDwY9X38cchmtndU3cEVDJbyNfuzcgXhEvh5GOFh233/FuqoMMUeNNGD
nd3lnk/mYidxCerxd3P9+cF1jOiB2fwdKFTZV5Ag9fkp4mO4Wa47prcpzywR7GmowqHplAVZ3XXg
ua0FoIqd2LvENn2IA2XsuYbwyAwcSukt1EAoYdwH9F9i2mDMQvjO9zM+rAxzcKkT2XhKct/g1azy
hdLa9Vg82NuDz2wxHjJf2nWPnH3XtqWqlRzLIcOGHdD57nhnfylZT4pEspq8XhDNFaXpsEks5yYx
6jz6vKx+lMURIypqzj5XZPVr3b5Y5CQQdSQzVvQsEfd+2ptqyYfqF/9LLmuA4ffRlNZeDejoVL5z
9sCnnp/y/cjcpeVduBqO/Ukrl7uPTGjvF06sOleMg5nsuNHjalj+iYoLRAYJc95wCUUJB5KTpYVg
Lz5/DHcEei6dVnjHM1adq/D51v28C3V6SToKIR30LlLnILdNMoPe5Jh8wHy+TYZUm2OgxAyht421
Zo5A4Sl2UCADUwW/EGASzjQRz7wRasnamH9QvjAZ71lodj+Mx9fz697uf+kDP1mBUROG6aw+inMA
3epd7M2Y3+t0auj7bWjYpM6Gy8fkjvMBHhgmQCoxCV5q3emD2GhWfj1YvvJKRdSrzeGX0+U7hJ5M
WosGqqVLQsn6K32FCOTQWLocHx9BjRtzamrkAoO8VUV0UYDJfA6OXkFSSakmPoqsTF13H5Q3Fa+t
2HqLJ4msq1XKH+ofojiCNl68k7vfAXsVMWWG6isXcVwZ3KGps8CZZ/aSJ+A0mA01fWO70N1RpjhK
JUkQY4darPACkPuW7xuR4xcOaxXoleifLpxx0TgFVsJ2RDA+TynqgYwo2l15gibhownq3j8lYjQd
5Wi4FrqZlx/0rF9aGnKnrwFADIMIqiEwl1i2f3FJFILzndq6bUE6EpHACGPOY5oqIgwaYqttFS7d
SIwry8N5mcFvXu6Af1N/YQAXYKma0hHPd5xhDlrrYRWbKcqK1NELmpe6RN7FNS9+2bL85NN4NJVl
Z21Ejd9DeMY4gVDFetF3Ao5oVxvbPnDOTNGtHVV+6vVQq3xZpw6QeUFZ+wSFOPiZc+6GIua9xJwl
E9daoe1ETIZaxo2crfO6FvgS4gJH7349+bAAX0nju5fSZMQvqMLAZ19S8cgub2JTwkpu/NiFY7ZV
NSP+LBG6aK5OrhxVKyx7PT28UFsnRKqnPwTW/kRyTrv0BS/ScIgMLJMsP5AWgOiA8/WEiva20sQG
9INSK9zJJd4GTCEFa/rU2v5QI+JqznZupXOJs8qOU3w9F5p4NTaG6q9E28uqba7GSDHNSiMQy2jq
GZzRnY8K7TYkNm7X+zDlIEQ3DYiVYTPIQYjQDHIixy2/UXoThqoRndMqwxcsyNfXXjL8B9wuG2xB
g12khsvqquUWq2I6inHk6Ogu1pvUsd0D2b830o3pwS2Sq9YYH1kC7RPEumwsrPlMclBocYhOxgpN
eT5dEUUcWfHTNTl07QVl4bBgHZMPMk0pd+2si8zgxEnk3I/lrE0CHIUmkvBLGaOaZjnuFNy7/XD/
Y+joSk3hni5p4nLdmEO7n8Qf31TbCmyw6qRu/lo9wW6KiDiHECJZ0PxnNnJtgTD0a4xiJ5BYWvOm
UzSMaq/zdBVyc8cQVjnCixcCNSXIui5o4CKHS17KvSgogT1oUStla0Po0b+Zj9jZMSsXtQEg1ipH
vCnz5cYJ1yxbxE9U6oIEuQ/GLoukK7S2jXrYlXZpCyPjlG82hA7i1WGDlHu3jZlQxIbqi9RcqV0w
1HzpHTPevQr5VGm8oX+zmlKyuJ3+HY3JM4WBoasYYt8fMhoL55+3kZGM10A2hHTOCPUqMYKGYznr
Sfb2YwR8Cxn2FuljPppQOmI6ohTJZbdCXwPbeumrj7moVavFHzCRxUiXLdCZOTOcAH2wEj6i4gU8
ZfDhLFM6nT5Pbw+7NBBVThDnOHzewSH3iQuwrxYiv5bxktRFIHQ/4hslV1oIasuK8KO9+hZHad0q
smY384HYscWmihEtd2scXjH95/2SGC++KDmR8HC3udMQfhu+tYe3Dlh5MfkYDE34Vdk16h2ZMuCE
2fWdnbfmYUEzvwxLp1unNtsQ5+s20Rw3J4Y33Lk34sD4dOweubZyKXOPXToclCBWJ8ZZ7Mrkggjr
RrQhWe4xsTL1Z+Fj9M6+8bQfzO8Bl7k1v1K+zckSwqABSBuwYLVzB7iMaKV5K+ZhN1Bat698/vod
8xeWIGU6s1sGAVHJ7plXuyUV30X7mrtI+jTKT01XtwSVF8O50P63Jf3Tx5P1ajPcy0suQveCc8EZ
W+2gzGONtVxVuMGGB7VG4D7azZSJ2tZyjo57LytJDEu4lPTvYZSXo6DDjm0EfNXjiNLeiTZ2rACD
pRbQ8BJRHjuESsWLObhXZYHEFGIiIn8rWqiZRUbhYE9qZ+vFExY8bRpzJJMCIEx+P7+N3uSuGQ/R
qP5hD3q4BOrwSggwd1IoxvkQHQn09tpxeJy9Y6STl1p00oit1gJ7FyESGdyf3ZRkAySEnPQzuU+8
HqK4Gde318LzcXnRhAxSFhl61zimeYe3uiJ8xIYM+eox2GAtrRi9pHiWq+SE5qzJixTnSKprGZZC
T/Zrz5/rMyP9BL8tHPRXDjRyA1ZyRrj4yxXV2su1e2Vcrku6cYNBXaJtvchfYPMmbgzEZBtK+Dmh
YTajCG0N8kgiQBkRLaxreB/tmjJ8+eQQ3yTrb1gMzZKgO/bpisbyZKnXar/cAKkTl7jQipoUQXD2
aGvMCfNK1stdDWURpVF+2lcbfRmO/F8NXZBvXBtSqO9mq5X4dalHjg2M5MRNjZxjfFKN8U5Pjj+p
1cb34IkzA7sm98+4QOQsI3c2ZKDnSUgwKTW5aa8KQet4lC2r9bE61YY/yqX48h1mtToCzm2sWa/d
ygu5oZAzC/cfB0cXJreDVhFWfttc2Si+ABEGuTrJyMoiH1gPgop85DhsucaZLxn3opFladMbjshX
E1Euc2q/F2LCwQUUDXJNlQrIsRAbZOWdOt/MHTdqby80x4VJB+6Xv8Qk9owCr6nNkbFw7dkb6ghy
MscnmCAFvUXL2bqaItEPAtwEOszHswhB8cKEGH1Gy1HiJy8DN3lznGxDypXT0uM8qdVBvMEX80kM
P1n7z/gqiEizfPzknltRPZoCVewj5NwUeNe25SFrkgPuG3jG8xt8Z4+kSJn+bFz0lycEMfCuemvu
5gNIngMqxJMojFmNShSZy58+S3z5uzGTTTL0l2Epug9K4AhdQqlj58thnKiKvIW3d7uLbq+AC+iN
mMGWCc1BVNqVoqZdOuhJxrHibZjJMvWgJxIHWZD2CBt4JxmGV9zo2RKZeUvaDS0sF3Sxn+CS9Cbv
+Vlfxu9e23VK5P0W6bV9NKbiY8y5Dv3GhkRLlyg0FFpucdq4/2jocPNRSRCZRFcXwj9HXZU1lFrm
VNzvSpAnU3O7K7t5GTALI6gX2HTcI19cIVd/FTH+wrYebo2CbDiF3HtBJvYprkd5zM5LG/s71zms
/WCqaWj+cGzbDNLPjsRWS7b0LZdtL5lfQ0NU7+Wvtu55m79ri/JHWn/N3/VInbpFEDPR5BcFxZpg
sykExQaqQvzq2b+4c+XYc3gfgx438tGGpk7f2+8wRVgE+NGoGv3/j9bg7Y9U/C+Bpn3l4uFrNS6j
bcflLgEFFwli7c1WuZAUC9HnSWnACDfbElN1oUr14Z39MtM3ila4+jQ6YN2ohCXLuLAjZ0gEgD2f
1BCbnKmfm9yNOW5gDECN919nEJvUbR2H1cmCAOUanYZGJQ4Yp7PCgfTL6/gW950+cLUqCiH6AxL+
BBpwec/k23zviWE81NlyY5IMS2OjLEGuPAH78WTWBMB9HQ3kkdbrJJwAV7cVwDzyMDo0rJawfG0J
rlR8PlEpjxt9k1W937BPXsyu81M1fIot7/FtIBcgU+i96i4lwoC6goM/jHawTgw7m5+Wl0aCfsOv
TFI+sucdpgtLPjWvO6+oul61cSjve8OUHIqi/Tjc/ZvFVQiRSK1OjkG0Iy/CvwHg9CfARpJqfPSF
YgkGGYr12C//bpoauSaiNBFLzx5KE71R8epjqIYPWakJILSb9zGBoxAa0+V65odffJulG3VafASt
Pf5zJE1Jhdh/h3f0n/LXkIDX6PMywdyh/kzPhoMjuaMQPP+yptgQOglhZS5oCB1AxaVcexs2ZmnS
kpAJtaBmQ803uOXdY7qjIR3YNRFVlkQZFqekIIyeTScI1p+Wacbk/jhZmaTeannobu3gvF3mRffx
0cLGOtK238jw5WLn77ajG1mYsVZh9UfJDe/BGtElX35H8COB27H5efqe0Zw2qKsuYXaX71w9iRcp
QQ6LjNo9DR1Cxv+YEP08rt63hFEqzEokMpaf3KaeoPbftAAPtfkNy4zqq80ob0UI/RWzv3y/7XbU
wUFPwgH/t0ptwQHkJqJomajgbhd8Yx5qv2LUg1YofxjHXayFzy2FwocJtCOQ1tgGh9KkaxVd2AQc
wG8lDPeLyfE7li5UuGTPXjL8i8nUG5Dwd62xKsFPlm25XJxLfMjsnwQPoOmBTqJAt/dh0/RcH0Hb
axB4NJYvX9SPbzsEi+DU3EnvhhWL9V2EAPsUs9cyqv98/4FdS2UAgSA8Ih38/OGrbyyPXkgDYd5f
WLsCbk94Qev7UURBiGkHM98nXKwBDYJbkw0voA6ay+C0aFYxMmw13LPrBFJP/8eM4ZsPvZkt1wPJ
e/fTZ9+M16AhMdjfgZDUJM4Hi/+XyjvwmV/By8ZQ+zM2FGPKf51PhCG6YObujlS47q+NQCsYqZnz
VunrjbAKfPB3XT6pmtPaTnFWP8NJuhMip0K1gLix90aLAJ8vJP2ztQ191ZKYjPwe7sd9TW/uxs7u
3kNyOH7hRfX/b6h2HlGXTLXGXoY1A1W8Wi0swSLni4JmcXKR7cbP75mbBp6jrn3NWYIahFfOXYgU
6yGXHaYbslnyEPWLfJFErhIS0ay32Fv3gS0wm5EmDMyxM6G2TWwah63S4+5wlDGOm5BmaYjOeDXZ
l44GhaN/OrgaYZ60HqUbg1HgukHErZ2NkgKEuP01wLSae2HEhl4tmM/HJTAGW8do+7OrHtHttvWr
8fcLPBejErXqrd1uGgV/J+dPr7ZEMJdQoi11Emuun/QRvwT2vr1np1I7jQeO8/LTYQGidI0kfSSq
hRy32h47wbr87jUwrQPHrg3FSFb5fTRFPceoUtubCe1Ha1oI7bQQ1sBudNqUsyW+ToJeS+RMcODc
J315r1GEMgYZdT8eakv7OEkco336oTCjOJeHJJQAUmcRdaXXD6zL7J2pa9VXtxB9mFanp1YZfet7
kug4IRPKb7Qg90m1nxHSA203lnboSHO2rz/zphZDke7ktzOBLgnjRnGzwubEhp7Hdo2qbPd+7hXH
6gsspgrg0/Rr085C4tDMQb97XZ6OJaYn7KPMU8yOj3Lu5OxuZDkLkg27G/394CO31/aLl1ZpSe2R
nR0vXYS+y5zVoKKftigB9+EkzFlD8dne1aqcN3bhu6upu2+rwm2FJkzNd9kRLMsTWSqICYDrLa2J
7EaCS7tJxAfWBjHjRwJveRTPZ53mJiPPO8cT2nRoNmjiLQ69P0gfA2G/O0ZZiO75NmA8AHGktZba
cO9W8Cgn+mBoRGLUdpYaPVbPXlJg7NZFwbNk6kgl2gYKBNo0uuVPtbq5l0lpdkvK85ZQbQxRHd7o
mKAhU24TgVyfv/X9V/+0gX5cdAp89mTd/U/K8j1DAv9tm6xS83iS7N4jOfEEqf7b4AmG206mIctM
6chtOZkLjsW7LVCkRxNCCyq2NR3OKaZEQ8vg8swJrMN8mIPZL8r2o+UXnwhWQB0T6ljAmI4lXY4i
z9c3AS1oW6tKRwQiyD6q/E7P9mrKGqCAcY6U8guUVbOyMRZ8srGf7yLzs/HjFdNBK7dHd7Nd5wms
9ul38fPCnJ1nzZ0/8C5ISyIJIxbuXzOeYvGfULTqaxtKUPWdgLwd6cEWCQAeAjSk/eG/Te0UiIzo
EVMJYbiud1NTBym76RYYx/0FAGFdTi7MRhPeg4E3yx3QVwk87ptczamWDWv/AYvzglFLZlMvLyKT
Wthsls8gwUBn8N1ZMBBiFJjX/dUzKK8br3chvuocH3xcA9HfdQmNTuKP5alOzvfso+2PVYH9kWZs
OFVIp7WN7sk5VQP9iZzsF7NZQpxtsqAMo2tiqr+Y7CrYk8FeQPPFhHNQQ2vm2S7mnenmAc3tvuqQ
t1WPILWXUEtgB2UukZff8Y+rEosUrbPUr0n18aswNojR5S+fpayxNyEn0PwA9sHCgYjjELqw33nG
MzUlfMBmLDbopxZP6CaSZ4Nxp/WroAw8LQQkq6UTsXR1GqXVEPyyetWOpaVHmPtHNvnGpPJzcYee
8ohEmLXuoNr7xuXCbPIdnd8Op/9IaRvVVIHKnvQzb7JRw2hV1NwdFXX2+NTycALMFl7GKxZhtCvW
LT2AmR+1gohdFn1EIKO4CNTrTWHduYOAshmLEq9N0c23i+FRHcvvZxd1wpDuQAOWqLmx55uroQk9
3Z4+Ao89KwfLJsQEdfMGtc/NhJjqW78Ydb+A+uyDDBaI8BLW1gr55wvoWst3oh376z0projiiB8V
U/21ofk36eyE/yzyKe+S6f113VLlj2upNND0rOVg7emByt8qZtaYPOZflVDX6UnuSVBCAFBezP4+
E1nwGXexj4FGv7bSv/Z4Wh5cQ2AFRiICZ2KJDPBjok/Gh+Zgx+eL82r2lBowz6S13G7106hkN6G6
pPJPbTjgR6h5zqjaF0saxjKcOMPGNSvR0sktuqE+oHF5zsMcHKWApDB8wStTXSUPKKNYjbDS0lui
Nl9JRbIrajKC6HjtnjG0S/KzPomYK4/XuM11SrlrYdNRq/fwycEIvqeT16l0o5kDe/dsp+29+gHu
Vb9ffjw84GRLayaAIXJcgmjlxWlUIOVQZmb8QXyLWx+LdtXEhQnSOKDP8PGnMb8LREKHHATjL65u
cnMqlXs/Kqatwi9pgLFdKdtWx2IGzXINhAn9+c5rqmWfmA+Tbainy54iKazGUYpDhci0OieBByiR
Ypro82OrJ2t50I2LswD/jGLPTVq3gyNFXFYCG+C6/pDRHuzaUNkNLTuSRwCTPMlV2vL1Yn+9vYPA
qmbiMyaAgO9f6QR/FWfAx14j6gBgpOTThGo+BTK4T0aDo21HjLE/s+T2uMb61a0xun8nwx5ooDXQ
rpMJAE/XLnEWFFWlfqwhUUjW/KU3M2/jyp4SOwDSdjdItSk3P2+UWBeVCuBFAQqf4kZJZnwe89xf
IHIrjsQxl0ALYad3I2LShrcTNPCr3/TlqjUXHexLfuN45cD2qFC/9RyR0qIdub6/7Tprzi31EyoQ
uen4d6TfcWwLc5YGopUAbJAMrVi/Q2JfR9s6G5/m8cOEanCaQ0Y11I+hMHNNLBGFImQ5nwsGZCcs
1QFu32G49R/k7jFD2Pf92AaP2plfcn4ygRsEzs0LLUTCFmoNjxgufv1Y6bjYBUDEEIXs1nhjAfr5
mWw9vGA9g0md2uGR+DUx/uTg3evErIGX1+fjHVZKTL7FQBmYx2GEsnRdpE9jG0n8QxGa7Xhbq+X2
bids3vU0IYu2cIzq55zRrGYRGtr5KVl/iYohsM2ogoN52kFBmm31WhDACfRGng5t4HAap+VPThdf
lJO1gbSXjVM+4ycsu+cACekgNTyY85oyPfbyqxnRoslS7Vr9uDptTHt9GxLcqbzE72xq5EfJf8Jt
HFagqi/1ZGDh3hG3oX3pKrpUUSM42YM0Z7lvmzyghqHLoLmJTYWh+XI8FpUxtyLofWjJ9SKCg57S
ELvi7xmYZ9lGZMpH5RycdIspnflZs9A1bvSh5TzMcnHMCA1YyqNKEjrYtbx+YO6sFgpI7EBfG3aK
96+Wyu2InN+nKSfD4UFwVv2rEpnjNA4SDsgT8bSCV2Ijw+hsFXpAQAGEUUA8omt6RQ5DIqdbmMP/
HRYVa5Gus3bq6UcBys+Blh25AvLuLsUh49MC7GfgA7riaH+YH253afemHqvOvn0OoeT0Kn9LE2MU
aqrJkCkmHNlEQAbktNvepcr/3GTKd/QHES4/IlvZAcJBVlLnPcNRY+58KEcjj5U+TUBXaJ814Zhn
c3J34fNvu8TsH9tjQfAvV/S3L8Zid5cPOw5X/MLcFUXMcUdAq1YkSnLLSUt/qI7l8PR1dPf1Cc0P
ZRH8aIiMRIXiZqddzLVUj7p9GC4rpTFrjf7pL23svzW2cwAVc/AhiWKHVA1B/EPHQI5wDMpsSu2B
Gxc4LipXh64tggsWgRqWBxiu6iT5LrzSCW6fdGS/AiHX7Sq/7IEo9Y9wN4EAmSng+AvLise2fyvp
OyNZ0xDp3XB1OJKSF8ErPPog6WTWlkkAmumSY1mEazVR0thUbaSID5qYq/6Jbu1HSjP8DmkE03wc
v6BsOaRvwZutFQHF1N+/TK+10tT2UO86u2s0J5ozOYiicYFzhs6ez0Ug/WzGlaIO2jfO7eXdZy2W
vocwYz1EvDp625TbqWAht0cGlEoOGYjw7Vt6863ufm5GFzyvnSAB4cZwVgMGDb49dW4zPLDQanKm
Sqm8JU7uEqctq058JVFAOBy51gDfFpKwsK6IfeWe9W67YESynzBIoKQTpiP31OROnmFFbWjAymM2
vNlP1GMulsbrw4Uj3NgnowJj795TH5wFxwZyYe5KTCbiBwXs6ldhb2tl5p1a4YGa50ovWcD7MWPA
Pczq6BUN/CUKeTFNLorS/iACsd36Fdf1xW3nXqRfNmcYN5Rbn8TwGVJII6IhAAuuewYdymhzAJd4
BqL5WbuS3HjtC4ycsKKui9emGISgNK/PeMSZWzpv38aLkSctGUEpGEJDM+9N9vvl0YD+sRBTVagM
9VrsW3aR6hjjeKHxx4ZNdcWptK9tpaSYM/M5to00xIZ4aXsNKqo3LwVmiP0uwdGEtU92EyDx/Br0
dVa6zz2VtKrUalOQwUfUQPaSpjsggsWkw1sUjkcGuri3WmeihM3XSk61TZezhk0CAlZOiPaHFJZ3
ERzEtp0hnnN5EbCGSndcAE9qLd9XnxvVZzSxxhlwzEde1ibgS4Svln4Eeu06GHLAvEVp6ntiaMHr
CB+ZdwY8Uf64/yNy+0YiGnTx0Uvaxxwe/JDQtVyduAbbxzA3AfNh96dUwYvZ5irBCFvdx88WQnbk
tBS5/Iy8NQwA1+O/p+XNsH8gR2ZSvBV7+dfRh1T5tQrCy8LXyP2zGi+SllnZgl/ySzsbu79y4+GK
XY8Zw7T/IRairgkP/PzagvBw9RiQtlC6IMOBTTIjevhQIglnsbYtLJHvHmldXw+SLJPp56V2uJdL
EdwIZtWl/DWIuSlCkEczKuJnsFW6+E2dSdiIWTHqWA63AdPgwPS5xq1oQxWVDi0q6Jv/JH3vCX9k
b67IiVpcuY0cXl3B0SLrIFcq4fcW4BhY+mxuiDou4akE3OhnYtXPLUmalVc4KiDfGEzUQqeU57bm
345AMMHXcVOR7sEAkmpB7vHgnUiIppFA7DFYBVl0/3WyfW8vTeKhi4Ouv+ubgmWKdJMdc+C65Ful
aAUr0vyXVjj35GRMdLS13cvO2WY+fFxvsMKwFI4kpefLTgQeshLdZfAuRmurB2DC11f4QSpm8TPb
707sxr4fSditA+zu7MwXfYog4P903KMzHxY5L9YrVrhvv6e5nLfWzwuIJPV9RsrtRt/Hgp05IjAj
NL0+2KJRcWvl0vWPGdk0DrR0kPN/yGvNCRFDlR13ff0Bj/vW3d9PujLg6/0e2WMEBLCvnOqMb+Q5
h+UILLpGYFzCMohigtJCVXNaGLimMDGEO+iH7yuwA78OY0wWVy/GDzl2hPjkCz0VboUQp48SQZ5E
mTONM5wWczr/DWlGKYKegnfQ6niUPain/Wy77GAZECwRn22S2zLsjSUvl/5r0/2vdAdIsFDmlVDB
fs7CawNkw43jslB0Di7G6TUpb53lm5F4CTxrEmOSLfw8rDzwOWHid+ugLxdaAlQTyH+FG5K3/KsC
Ba02po7Q3ZVs9HFxsir2dK896006Pv3bgHxODBkJ99k0jb1TDzxVbliaLGu9LH6t8PsS2ojHIDx0
o+ZTonb1mXdOc/0EsliAnmBVcJYreNvxn+8BWaKxzkDfdqzZWKGfX5g4OmoQqJHKSiIGj4Qq6zPI
t/SV/pIWH4IvB8jU1w7ExjAW41VgNg3BqXs61rUN5tbUIGVcVLsz5TmQ9En9X8AXgA/JKQVf73JB
jO5SFXGgs+w29PECaaNP5b3luH3zhEggjqXAt/pRPq8Zt5WtR7Ot09ed4k7eRBjAm3A2OtCSWnB0
MxcSCZWOd3DC2TtIYesGjvq7HztSp1ECIzv7j2qpaMPL9bVB+H+SoAExBmgYlnDXw7clpIIQEAQO
68nyP5JL9rUZ4dCpwf48kx6TeAioVri6ycC02CD3TCF6FdldRE+dVWTKmUFSNb0Lk27czQd2/BJU
WkyPhL8yBsLCiG1ocYlDoW585K935wm6PWQGLzkLNKTsizynn81lUoWf+ecX5Oa2PAyzU4yDXZMn
wuklmGR+KOJKpeRYuM4Xva5p3iGG6v3c8YChKEWm7MW9gqGleNMahQ2QmToPyZMFbC6/Y3a5gSeF
UBWU8RaDY5t/3RORdkQcwaboQRM7WYJVc3SJM09maab+td3DEnBVvCvOwaL8Su+wVCe9A4kofmiD
tJNzjOsfgAaQEKaNRJlytBL1aTmue/GNpQ/S/2+4b94scY8QRYwerb+vPLdorTVmzCCSWd9O0h58
uxARP09Vsg35X0ofmZrWwmxaimI+K8a0SngQpRlpNjA7k168wmRodB8wE0gqucGqh3WWIvFP9oHt
K35VmWWPNIJJcxf3uMSm+/jJRWxVUBx9+2mdAJMcaGerlwu0w14i2zK8cGiMiiU8H5WWcMb24wB8
Gsd4JfnV+nY8KhagoHFzw45QhwuvK5nNCj9s7OEtGOYYxz1byRPj5bKx46273vQIMm6Dwm3VS8mf
CBslbr7nkjrzjXq8VB/KwkZlF3zMqoFUCJKgr9dKhEfm5qpC36GvYk8mPASufCvN+zOkX+93rmyu
vlLn3RuvaQErTx5UN1I6vV9cU065A6BHVS3F+RUaV7/avV6b08GxiDuRCf4l0kFPS1/7SL5GvrIf
YCXoJf808dxIHkgyDkkcIctmgpkxanvKsj3TkSQxwvZFJsQN960GSWxXDz61HoA5ylo2yfVJT6pz
JszJykRN5wooldyqejE8aELK8guKo4cGr3AM+kwM40Ogu9lUChmLsoKyoQeyIOHclNRWt+B7ISfZ
0EuyuTKadeTXr/QSenxYtCaQSJQVpimZ2/xfVe/Bo0oD4IqTYtvVfSQaUCi6A2wbxy1XrJHhW46p
+j0ZndNB10YgYUFmXjLt/btXTCgDu9E0LTaNIgn4X7fUUCLICkCxTXG+6jtCVcS7t3Sz5UYBNw2I
DKaq3yAwR0zNHPZ5McTdsJ84QgE7xhcz/S0/9wjjFW6CTvmTAkU+LEjsoHf4CmoaZRvaJopfmghf
c3/4PniM0XUaaYLc19+yF+d5uelNaTvsHFQXvCeQE+hqUyr/qkZrWCaM83JHRigWYebo+LZqgPPq
b2L5TieEfGjNqQeonQdIcch5PIeFmX4M4TB9xw9DJi5g3tBAK5DcCEQzC65cOSFms/e3GLiBOvQ/
k0IzUNw5rbowSgz/rMtv+iABrEa5jzMKY3lgCFvZgWa004DFWRsYvS1K9lOzGK2BCAcLJ2+MI6lB
HVqxXMkRhHBbUH0+I8jKDunopiGGq1P70mym+m3QKCnRNhJAzrTJ+eIcXn1C2hYczocS+AtONxfe
UvIvxyWIhIf2f6XapAt0g/lfjyFaB+oKd8YFxHo1N7MBOv0W9f5KTZh1egQCutQwhHM1VVVbQTYV
4lkoRVXw8mGe5mZlQo1hDk7clMKtMlMg2ry8SQqlW+RN3mGpb9MFGmmLjnqcbODFLHkBtKKaTIvN
KLslRqIvm2HgNRfaCxgqxAq+Jgzr52EJXLFfYnOP/w/YDvlsfi5/nO+RTsVQwwYHvzXCHoI8ITyQ
reFWVmyl7qknWQtex9BBOPJdPMYg2ANWxN2YrT/c49LI77LDBOs6a5fz2eaB3gnAtp/6kH9RFxiP
9GCR7X+fqwHfMGXhqNsm57ahF/9MTAipLw3dpNZ15roIwLZyO4TWracfbEwnBFnf+ijC3QqK1QhL
p4gtI1+087JapZccFasZS3t/Hx1HetencNTjM7zmqp10eSv7Vcre4xNxtCr7kuveNyJn/5bhohGh
PAFrX0IZW6S0pJIwe0P0pyH9vIobn/IuDFZsnsizn4fJIt+iy82J8IOdacK7OtANez4RYJ3l3MvB
oH2d5a6JDg76l+eVpoPplFqVJporwnqUblBD9ZGmHbp0n4jDkyM/QjA9hnQofuslLU9jFjJpy8F0
rt4k283HZ4FEbaUkIkKk8DZmaieLtsGNF2AdriEISvhX8FEOagTwe7j/O6hSApJ0/qpXNc0AgQPE
Mnp3Rh+E1XfJ+20F17wcEsYeVHtFWr+JL0f9S7w4IuZayjv4+ECTuJPtdi+x0vmIoiMcgcrylIQ+
cJkwcNOwM6vqzrgN3k3I8009RE0Yv9W4GOZDi7qgCf6+PbrowRDGR3ibOcbbA+Xm1Z3wUED48XDT
1KwRiggyzjCNFI+XUaJjMFCLu+ef7fAuTKgECtQJQOz+XrsIidBpTo5Z2lT0k9HdE8ak8xOOkTpD
tYF4GmAGIc3ul1E54QypP6t76limyC6b2i3ZmmlfRJ72CLiXJR9WThrZDkulgbKmphjNZMClCDOP
hsukxRtEHbbJ2mOOEw+GtoxEEQ4S8J1qRVHiu4gtak0HOolMoz+EQZ9LV7RpvFaSZden2puZjGEf
NGBk+oH227RsLQ3m57n1ehWDyRQK9Lh1P25Iv2Jj1j86oy5M8Iamg+Qxqn6LCXsT04tMVm/5/qOq
8jaOcYYCditwkZ/45vSPGxJ4HoRnWRawVC/Z/9SHhf+bEXIssxUkeQj1EPkKT0QQNS3uddfur1ON
IP08R6rwx8sCpDxQRjhEjOU/4UjB8HsD0JSiwihgW2Z5ZNYFfchtihdf1fo7tMEKhDVfVJ8sd0HI
D0PHt4UpsDWez2OS+HIdTpyfRvbn0zEr5QlfO6kgOihY0jT9iHPzrCm+jn2xj8+5lfUWCNo6p9bx
9dhK9++mkfv3d5cGZda4peltjtVTmCNwP6WkMNgD8lxF+GvJCln2xs+zRDB1vjMMtO1Z3eB1RX2j
oEHHIYjLvOrlxJigfOSkqBnrkZMTweGGuoWeHVWnQpfmuw7jnqhUiA/xpOID9FnL9SZAFqHRZDF8
EztLiDQv2tbpkWccVww9ww/VFR23J7OmqMMcTbK4YcxVXXwARRsllnrMFBd4xaPHYeh5TN2eJ+bU
KtDniDrmHYV7w6WYjHwlHigP2GvcjFvU72ksTOpAhu5RlIeMhGUycZFIAEkVJCNUAlfRwOXXwyE/
cX7s9my9q895hMdezJ94nzLOsetQzD8lJdFcmy5d3Hp47uw8Dqj1sckCFk737a4R0YA1p/AWDxK3
WzGI/OwQruTKOHzUyVPqak1yGMxo4MVz6slEeZWr/JfboQJrUigJfIKPiM9nsZ9zNeoLFZeIknPO
C42zEur8/MosVIPRQHxhutDEjW430BUVp3GejLOvDZCJI7m2gTMWmr2jRMrFYrKmz0uIqrucC8WM
V8A8uNFEZUaySq2pPK6OrIFMeyZUEZtsE+A6qrl4oEbJdx3+JAWq7OR8+qgAQKq6VIkq0OkkjwTa
jAj96e1oGFLozKJjkqmV6lYyyGGLCMlWK3lz5qp+7s32rirw1RpJRd99kjogaye7yOidRZGw6O7r
i2OfNmxpGJIQSNcD359ubuuDzR32orErQzSSRvJDJkFe+0dfQIWOug/bTwVNARzbt67c4m2M90J8
XZqKW0YYmMh1chBwVcXOjmmhogvfSXuNFhglgPR6t+OaxqgS0YBRTkdwb3NrncSGB1x/t7Ligk9w
VZxkVY3BsADN7rOLiW7OvYbPsKrTYtAYBfj6iPGiFPP6O58Jso8QnTrFbghsae7bxP6/OBJDfYlt
BtUd3f6OHutBGHwpRuXI4G6Rz61AX4+swG4mpoMi4HZubNA6eHw8Uyjt54crevFTmhup/PbbH7NH
rZvZXh1BRqlyCp3+9O/LQzlxb7UNJ1Z8BxLcmMLT/mYvr4tWrEd1ZUsmjLM6zg5CdLBCrCCIRuFL
zuAF29FD3hYU9drnWKCU4fCfYeKbcv7j4yG9nA6v3ha3g1MyegQupvfvAC3oN2psA/Rw+hb9TQWA
jXteHGVB7EzecKPVelqjAFIUFB5aKPPj3tEZRYmB1930BgCXotw7YM6xrGmBYY9nJnfkNskTRyVE
etKCliGkiU2Ce8buGLRfuGyv6wcp1raUaJkNfX191SdZM2NN2e2X+NXA7tLr++1EP/KwWD5e9YW/
8ETp3h7qVvKE1ldowG8i5nQ5rvVsHi6PvMfUCRMfwh+Le2W4IU5xCkwPBwtE/P8CzjHjWNFxb5Uk
eKRNylWMMyWchg34Vn6l
`protect end_protected
