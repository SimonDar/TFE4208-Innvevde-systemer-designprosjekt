-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XM36QnuaQHT8GbQGF5a3FYi/BXPPsuMll4rTjyXxugPWcI+UMSwpgNcZbb+xTnZvVxyc1+Ngc8mC
DXvbr0icOH737L7Rip0NkTQGQwCL+Yq/fRW07NzXDOYgrp8IniutNK3I5blNfOoE2mO1Yw2H6A8j
1RTcPAGdj38K51YWxqROm4uZKR04KYMZ5x5VLtOFYiKtIXP8IB2C/GSXEG74UomC0dAzhV8TXTlh
BoNQjO6mWzP7wwUB5i9qshbcTgUTORuRqUjYtocy7vZaoI+h9PRDK9pjICSItF+bjGK2V8t5gtE+
cFpGvLS3oW+1jeM9v20DOZu7Dc7gfXQ7MgGeQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
W+cVvsmN7v88Uht++4YaL/pRDXSlOnu1BqzOwBOOkAAkBZx/VFKyMaS0x6DRKin8PHACekHMzYos
uJE8wCJaQ8HVeIIWhaBdBe6G13wdF4dY2VJqu5IinHRCvaLhlDa7u1QqY0AL7hLwtau2WOrLxxYO
ox5s9DKhFNIbTSBNAQpXD08VmEAOprEuO12KTcFy+OqVE+HOJ2+fgRPUBkXRwffp+xlh0/bjUBkn
ywrmx4zNIyTzLyD0DyAXKGkOQiHIu3ckwe2DBAJX8vmGjcBIWviUIY3RbIOsp8sjN7LBVME7o2tH
dBDwUkPrcOKiV+1ZkakQqs+xGnRqgjpaA2uJSDqNHDCvP2Ln41NCQe/VB+fb0eimLiKUJttRcosE
a+utAnZIuwrdhKEn+8Qvee1L0AvimssBsX3KO0n+PYk/7hLVALaUfGfVwG2gAVG1fPRARr6a1sUk
LP1TC/yNdbTGmykXzmXWHewfEgHzq+TXRRMiM/wkZ+h0qW1BdXMzmPCwMsQkLWqz+Tq4gR44rEKn
JxDe8laRFMd7xHGJXGUHgcD/t7+xG/CZvDKeMk3RQXVY4XOTXyndg9eA9sQI1UuSNyOUEBBTTpMh
zH+ZeFFa00H1JUqzzDwsCw9/zRPVhVLq0BgUY2AqbGfMfy/57l4ziugXFBEQ6bv4J8mQyzu2wxJg
gaotIhG754ptFcn+rgcNFP/xBUaap7x4Ary6UApxZ/cqB9ai0blyLv9zGGTVgYSap+a1t7sBIVYb
8O1vUATQTNCOE48mnkXZkMXVHkNwcDVLjVthGScHWGY72g9d9oUtKCneedMIeoLimqfofF80EhmL
8rAefTMjyLuFafJMN7yXRZhCb2Ve1/o0pbT8Ex0d04v4MD9TCwAHu3s345TCdWPdyNQ9M/jMHt4Z
00/Ee2L8KFVLfc2o4bGh/6lo6QPqeV/KHvRiYoaAPs7wZ05D+4rg+Le+myY+Yj4WlfwSdg3mFoqo
HlxPeBxB5Ew+NXoLKMBxL4Ldmb3fOapqZyzvCQvl7UbYeUa33v21jeYXtzK/fbbbk413pMR0xKGF
Ibcu7I4oXasCPOhVmGvTiXcy/Lg2H9QCqhqJNiR85RmN0ChwlGI204ZHRQ8FV8mrjC0NIlZf+egL
Oou5PChvWtqlhWRE9vKGswu28IzZqtuyrSV8b5hiFG4AJnDYCJy+yS5LTRCt7GrJrZceCUndvQWG
Ktk4a6AxnzQmuWVTH9dJKZWh+gE/WDCbGJwCem9Bdx8rP5YYZhjGKS3t717M6o8CmDMZ5Z8BNm7/
fFryAVKQspQ0adRkASRQIluT2POBcmFjkHKqn73EL0752TR9LVmfEuvt7cy4N5NYkYj+K8abTn3M
SGvM7CTMZgDO6kDBHOvdf38g/Xdr7EHcuLpB0/kjZ2w5F8bIMA3bGu2vO8ylnM9NmNMSqeowvAXq
1wX9fTt85YiQ+MY13tvpCBl1hJ8GAnFLg7ReFyLfuJrzZk2gicZaCR5NRqMTNpt9Ao4IAu/QrHd0
m3apqJN+5P0APiC5MpNiZv+kdvt3C8zCJmw4E0GSIg75OLLnr/fUMDKskD6qIVcu/zUtEeNETQP7
BAmmHykbtTzURG+Pnb+p3gGX+WFMw0EGSwBTZPQbRWzcKS34/GIuQalhHXQfInqKfYSwZsfJYhzY
/H/aqIFJ+cVg+Vsw0M1Z0ZMlqX9zB9iH7J4eTd9tGLsYx/HzDIYiR+xzohAXWJiYeGLdGtIXuXz+
/+Fx0SypZkIJb1u78jk6i8u8bFebldMWfI2qcSZJa+5JkTa+sipfIjX+CNyvvzEBlwcj3TwRHx/3
7c9KwkG8kzeqHIpBEi2WI8e54TRQuRha1qbKO0I8Qpd8E3EyUo/aliQUAxG6S5z6hH1cnJTY3cdu
4ikwWd5cqlEUQKJZ8ZGRTs9IlR72Zn3qi7X8PQhp7+3IXRQnPIernev4OoT91ud57gdgciAKvVPr
zBvzLXk3LAclky84j340ETQ5ni8mrHsbX3y43FmpJvaFl6z8GlawENqvo7jtrwWWDZytif5VC+9v
YH6q0qX+3yoTkMVEcQ7ErHfC9TxHm7ryfKBW12oHb/Er891nOXfjtUUUZGN3HewzaLfhjzYasUvl
bmOZ2crM/hbp7gk4LzV4fjBk+9q9DnfXI4KZDTa8GpZolaepZU/4uzW0CLm9ok7x/HWRB6RTiB1n
G0ipkgzy5goeocsjeJuRI5aj8JqH8bKiPSqQ7fvyQ6mMp35Ldvitu3a+veEmgrqFKAWz0eM4S8Bi
ON/qJ3Bt3LoRgYUV5Ym+nyWYap9OxPNWZ4jz0NY3xhyz1eP3GJE4OI3Q4rFMn+P+40cPi2ZiZCXv
owYGdCtoGMTnQsfEdRik6LGQDBTvgk+Mo8HYd9xyHQL3rq9ET1BkMFSj27a66np6QDQbh5HH5WCT
WnzHYH56VImWauFKcUcWKIX8YC0qZKjmCer2jEEFqgQSD3+f5XTpe6N+My5SYVzQuIlzVpwUHtaO
jAfzFzuZ04hDLY9wJNLPDUmV7QXZBNYeDvVrYkyZc69sNrVnA2pbn9zWM3FQq/neakmFtLfsAC3t
FsolmgBT9gf/jKcq4fptllhgQJl+mtm/HRz1EMymdlxHkH2qvCaQOqJwrLPATGbqAdmjyJwoH0be
jqnkEB0xzBqd3J/Lo09edB5ACC/LASuhTTTkAWmCNOEDL25kaE13NJxSlwE6101NtXNjy4wAkiit
jrUunbDPvUsFQjr8UBSDPz9rYP6b3kopz0YsMgjN2TII0vHHaCsFYgqq+4Io7T2DB1cFkhwWxuaE
uXax5b7KgejIaJ1dPKtQhRzcjSHZlxpftOKk1yd2LESkJACykCTxGIBIZO1g5aKGPu0eqniAbw4m
O5WVrqC87oebdYqxZIgytktNeI8Dmu5dCmH862iUFc8t+1mZX3LdHdr33VAV0M0+zuEWsgyO8xHk
YlbtuFklepxDxmj/l7iJ7MOEuUHd2RgamlOP9Ohr5xGfI6Ja2Hl5ptlPNfDsr3GX9iTtSJIThwhR
re9FuQeR4IcLLfinfEzdGLS6pYcA3k1Xmd1cJDWaw/VsOynj2175sVf3PJ89ac7xCri/Oxw+YPYz
ELa+dvcw5++omqyfVAO3GUtPqn4+B2ogvmwtkZgtcEi9UziCq1nvduk1M/CHU5mKtaxpgJmk6Ham
3Z0i+htpqgq+62+1H5p1BKSuQV9YmetLo896jRAYgmlCjaUEKu6IJRQYlGNWl/V+zkxYjnUxfvPi
495Es2kjb1lK+TisNigCfVCTXPp+5FIKR6srUX4x/C77cjvY9D6CmAGJHZzUlQ2jH/21b+GKMl9z
c3FbGd4QNtSn13uXtXgwcgSHwb26XvtJMpgXTS1MLd0FSRBsk1hzl+4fapSKA+u7oiz8jrQrXS5K
AjFMSqRfx+znAd1KzTTLAKuOqPS9Tc/pCi+TePZi0tLge+KNHRYHuOQkJV+xakVhaMk9X03bcvZ0
gK76YkONWj5OBCe1/OK4NL5x7fd7Qx48JLLSG65G+wHN83nlOnlY+Z3Ccdr08lLxGxCW0p3ZwdrK
Eg17fPRDr23uJczt2mARumoXORxh0SGiyKOoFLF3uRgiglV4/BJkUs1e45HwX+UlHLmBmcbD4+m+
Y0kQS9WsuiN+sKdXHvMpnvVJwqtp6e1DXXmI/P2nNJAUmUK1Z6AZbO4tmgyEuuKgsVMREw9KdWgU
o8kSvJxh4PWKTE4npnMQ52t91787STJm/Sjl0oP6ZyeLRiV1XrFUwWngz5c3dSkxkFEcYNz7ohWo
Hcz07UKf4pFvHnKKOE8vXT4WHcTcdAKJ5LdfeZNCuSBL/VGA39IgwyfTOl/g8lXmHyiUPvPN/8+5
zJP/lMRv4q+UJko6iM37RBFVxmkCqvLS43Kpx/SAgPwy/X5uoMYM73xnDBBCdNhrbf9kKTSaHVFf
/JoGhyEFXt6fz/AxXra/UoOZlw/x8xpWnPXF1bBzyuZULssvivj7pG1pYg8srL4DjqOC37PS29ZE
YXSufHQbpRlWASj3k25w77dgHIXvWsJsB5ZtW5rsl/HtMd/4J49jVUMO+LXVilRVG83EWFcxqgWw
Mu2VkVadssqXKG6vOhIk2JZqdXRgFrU5fS5I6aOIohevXRT56BCMkzpEpKcLt8vDFRL/Yc0Fz0a+
OCpiXsEG7byqD2Wf5CtOFceHZGvDHV9ozf4XQTlO65bMxAiGXDDDyMQ0P6Mh54VGnZmiuC0bzp4R
ihIPXSVWmwHCtha8VaarPKU7UHiCl33e0Evu5C5NstoaO6iYDnBFdxwcSHY1Be03G3OmdFToUep7
JR/mLxXO+TcMnc36CAlsjxx6p9IkPtJKuF1lggVAg2oNTi8Ftunuv11rdWpVnRNrmR7JOiO656QE
NXQ/7gGJb9BTjREj/LytpToeCS2FCk3pL03pn1ZJQSdaHl3pcLOSvp3pYh3ErsdJMG2fNHnTb+ac
sbWpxft4Zl+meWiAPaJWEvw5HciBq6NRqcGWIw7/8oiDj8M0odv4qb+BX9DmU/UYJ2R8gHeAEl2D
BdjB5lZLuyJhkXF+iHVQe74ARq6LkYw3PzLW8A7iiS2LL+oXvjbgDKUztGcH0jL+m2OtKGlEY+Pl
gCmLvAWpDH1h91x47WLddDIY/g3VavZBM5fE2Zaqa/UZ7F/RmQldUe1uCiY4PFJIamQGa23oKy40
vGiVMoDFDRWkGdFgjnGz2rRsH4a1wKZYlHtTj7aIbTgdlDzSoOxwQdTFOOGmtgA2dQb8WzzawHzt
aSHSVDSEOLjRmS3FToXA/Y0Mh2M7R7ThHJVJ3AKfJQl/EOyoYLiOdohg/lL3wCjXCkANc6JHzf0+
9IZcB+Vs8adV2Arzs3dnWOT7xz6rBXS0gpk3WEU1vSpxvBG3jhaT+EJXQe8+YV+Rd/Sv6roozmZu
jBO99jtj9Sc+JlOo5FQYZUIbE1EeMDu4bDruy3BofMk0Ijp4VKlXbztLSfDW5IQuetgt73XYc3EA
/PSmdIQyUPNKXwiurqeKvwdceEhTNyWbAlmGMYQ2BuQKitgzm/T+SKAXLNN4FkwQQGON8Q251JJ8
ZM/PIUkYDO7L53k0g8y9jtOqXzFuP2nP5I3abhRhWnXq0X/e4CAdcQbIWy+oZJYowGijSgC6nl2y
7+7kEYAkJmhTq9NkNoGfHvYhWWVMRbuaqCnk4Vb0L3mm+YvsvCopO0fdQuJySa4hVyE9LS/O8NIM
sh+ceTcfGks3UsYVVlIfy7j/Jm94ghppHpAvwXfbeQOV/8hkgcwKrjEK4tBbB0WtdqJb/5iQ/Y3D
zeQV8rg/QPBnOQ1iwYmmoQuy5irVsNDisTZ8a29SKE+jRNA1+Yp5L5tMGFvZ4tTipcxgLO12eCON
RsG3SB91fRFOXpcpjZ6sXqtqGHCPCsxPbcIjhxMFcBtTdOhUXf7ZEZPs4qVf5bT5YDw4GI9C/jy4
qd9wm06YJdE5jIP5hYQIczlsFoAEooiKO0lr4L7/asm9QWuzlE2hmncH5cGA2+9U2VgesSIY3DjO
VWhavCVLTeqLJwGngPyCK37RFdveCjGEUduJTLHG2DW3DWDhFsW2aKD5nII3z/qamOOXe7gWd3e9
o7ogNrHPFHxfWz0eG3cfKL9XgthtpUw2rDbROEUzLDQb+WXyREMPQCsYlUIvzyL5AplbnndJj3w9
ZqyK/Sf5kVbUv0ESLDf897wi4qoVpeJ4I/wzr8onHFOFv1lLGkhOMY8Ly7GGsE/fDODhM1pwsIqs
NlRnxSdP2+hM7wIdn3IQCrE9Mse7YOBl0A2HdgYex5ftWX4wVZaOYbBrsANqy66fQz2BE/CQR9Wv
OszvldEmEwmyhq90t33JHypQuTXwFgUX+6+pM28I3RNLmJmXhs61AqptK6kshlVdCeCHs7EwV2bq
8WQw4tSvpqMBszsy4Mjsthp+/I1Je5Py7kOHVsTiP5itVi14zonSuR0X/SxfXH3nOc/vPlzko9wT
TLbpn56Rkb/N1Zl+pwbr9bky3jZOFjHlg+XlB9sQWBxfixV+BhcTP6qUwlh0nZncdIjz16GwS4B9
PWI6/p1LDnCZ1snDxAhmiiSM6mDLcoe4QEcp+v2nEuwFFfV+OFU20pnLW7KT+YKS+YVKg6kBLf9x
5DU89GdDkoPTnBwzqWJjct6jt7xNEaLymOUgP0L0WxZQLxiOE7zfWW/tlq5AHvOORFcQYXFML5y+
0HuNioLflRM52W5Fx344fTZChOuYJmxXuJ5COcp6ZYd69bGdhAXRpehvZawflhiWJiFIQQZ8Pe2/
N3rFBml5XLscMuhzI/31JVXglEO142zQeH83RbxfJ6znYSF7A1wlRyFR0Sg2SoaCDcpLWINZLCfU
j5G126tWdiUpTfZ64j23Syurqz3X9cNe4SPyltvXLc6R/UCFY4a4CDao19ib5O1VfYwhYbxHk8oi
YzUoVHLI3hFPn1q6n4dEfcwNeA2icyek9ZGUoIfILZQr0MAPHWbKFGQk8HuwfbY04lzd6wuaWVai
obx2o5VZEDRf6qPlR7+kEk1KbTY2u+IXJ1gUhiDQ4SUYs9BcLxNki+iNnT2oYYRU/C1xSjYeW0ZH
DybU7xnvTpidA+F2CTgbf1JBTknd7b3MhpAj/iQBpKDY26Ys6IPJWwaDz7SAJNDOQG/m7/3EV34G
FeFOQLdWGdZv2d9jZuWlcNQZmvJvCOQnVdKjm5oVQxwEf/W9MmKynC1ERhPY8KczZIaCRGATi7l0
5Yv6S3VKRXIoPosvOnyODI/8wOWc0SV1Sfs1SLree5gJhB24L67tT6Zw7bnWzKQcxTM5kwMN2rvw
Ds6dGyPySiOOibUOgmTW+MmvTiGfbXbGXnqYxIM+E42s9pRIYlQ5ivRZIN7o9LS3mq5alE0Kehrz
57wWE2dkDYbYn3xU9dTS5nbQ6Fw4hwJ97jkLBpuZC2tOQodMlPCx062eJsL3w9/AjKMs8hWL8aSI
2C0kiEBgKXNGlZ+JZ56taR/xvDLqo/aUZMZoYzgZZIAvbnlXBgaOfiPlBimzQaP7pcpgBj2vAl0u
oa4DI66OqdrqYPPmIk+FEhda1Du9kCtey39aIMaoak5QxdkSNEnhm+oBreHdHqMNKMgnojFah07Z
Gqa+jUqsiKTxdSihvGVop6RrWCOx5zwOAjZsKATMuECxbx2851bX7fPnwcsk1GOxDLd7alIhttz9
U2+pA6wJ/F02DNeS5mxIHA85jT9Wxnnp40LmhA/fEKHqS+ZK7UJDiTIzS9jCxZSMsW3lTMJBXfNt
QZ1ci7W69tssr69K1KTAEKBHUNWBA2co+x98Od/y1jxaJDbilCZZWlnoplEA0FbaoKy3RKgkr9pt
G7mmzKBDxZ/AbwrsjXy6XSlmbflbYDy1M4rAsJOoWcV3aY6eNJ9G/76iVGQmnXUaeXVO0SXlDCXg
IW9SBK5XsbCUf0i2mN4wkfjsbC7+WS8nc5KMU78IgyGDkXnl1MJbz8mae7FBTCMbtLWZ73Elg8c0
kLAWXeEfVoxH3oS47ar6rkkcczLQREWwZJYY29D4WS6hnlC3ewNGc89RBz6zVXHZrrB9oD6XAqOK
ZMzazzQm1rm9Iq/OVdO0AE2gAP+usgoKM2b+8nMaeZUWceoVwKgR1K8qJ5oPEiUhrCY9i8VifUEh
iLGxl8lHd5Q4AEPZYaXANzbZZL8WhX97A62s0VCUvvjzNeIO5tBg48Z+SRi/cewP/Ytx1Ajbn2z9
N1Q8aV4g4lBgBjImxTKrDPAu60SPEbgif1eGkSnZcz6Tp7z76iBK95KWzgtiVgvS7NCZgimCe6l3
kLoFWDxewf5CaAZK5hrwneZ16aFJAf5twVCch6twgFQYZAGdY8C0q/J0eb2HHvU3jRwpHK7oKBqv
mgwQgsXzjVU2mLzaYJALS1Z+yFsGGxP7Gy+bL00ZrfSrtcjBnBi5R8QAi2KKcJuONkxO23wdiBUe
yb0bnGcCpr6eB/r7kKcis0xr/UOfUsvinrvtBS8YY2tu3Z2uC/tMDhFJ4RBF8wbj5jyJLbGELhAN
i9p34OTSBeHcF3lKuce+FBYt5eyN48Yix1FX20tzeLRCdE2z29V071lv+ifPLvUXzfuIZVWxnhB8
s3MSlMwQ8twi7D8biG1Q1gv+cEcR51jjcE+1gqZzQpyFF9N9hdXiwJbQUeQwLbjZUjexmGWCHKOp
4JPusjZAJVGx0uloW8cTlW+2G2GKh8BbIa9G6DdOCc9+OQ7/8BhdoOVylNxbnueWoB5hZYKyv/bA
tB465HCRWmW2D/r5Un7kgg+Sul/lcEzAQlghUGB5qlTLbNnV61nUsLcqsb/lxJsG7FYz+5PTbfxq
XDU6MyQI94gUinA35Z7L9zaccNHcV0gYD9qtFDjakIj2E8wQD8uVwMcNz/nlmt7+sBIvV5KAnW27
PaU8uWSSHqRdpOkuP3WGES9lF+5I34H6qCYZzc9gNyA8KVDyjPrFGnLrEJdPWnUKwN/l822Xn2kl
W2KTChHXtKOID9TvXB2zNdReYnTEHQRiYg22J5p/T1AI6ajBtJ78ndLLwFV8WUo3InuSjChkzqJL
1pAHrcIcsw9TIyCAhWksInNW23yv8Q5TwYFUGLrRikh1Dwk8MDh4PDnAZG0ar1AA+jwenx+tf2zt
L3YKRk4TjOoWDSLV7UdhddvnioIPGvLWCfHIhevv1TWaxDbYgLhzP9v0RViVC37ske/ghb8JgTko
h3hy7TC/8iXc4u1RuYIK0pxwKzUOXutGMqOIpPOWTNMoNdiYzahxZBIKY8ZsxGMdS7FnAYriL3wj
4fNNtGgC6SDF/3/i02TY6IYOIQzd6sCZM0wCcnAtFjDvVNGzETKdBHTJD/G47NYNEikkTMtJi3JA
tuv7dTCLyr6fg4n9adh1AjWBx/1XQC9PPNpeKBobhNrSgRkwM/BZqT9R5A9jS8+cYLtXu+4SHxv+
JnwAIN2vPAn6iy4A79acZNXedtt+cyKOM7+Z+exBEQ8RYqfLpp9Kt6EEo9ZuykMXkOIGRhcMgqa9
PvbvrR6dRPdmk2H4K4WHA0mnS+JWQEemZrn3LjlSAHAlSILCVpGnWsa9kWKffR2VgUsw0hI9rX6D
sobDGe5lOv/4bmcOVdldy5BHtMct7/P53wVw/Pe7JwIQcmX4FX2wEAffQ4vG9xJ81DQgt4Ef+6Nv
56z5WzQzlXrSW3zOqBMrKb0DCns7YK1RAOKVaeBU1zu+o1w95T4r4icFrebTLXKhsT8x2fG8l9z2
GNqcMHXPvRLNNLdo231n+K9Fb+FqfViGA4oKV3s5rkHpplerLtKyFadbxO2S7N+7wn9aEjNwkWWm
lp9ku+fRVxiVf8N5cY7zRJLfaggeXMtksQhpJm0ZRiEmP/fEDhYgsFrdWj+TV0Lyg99EZrlsP/Nz
OjZq/d9/ZWK/ckJ8ybZIifpeF7vE+6xaJuLq8DViw4pFhwXEW7nTr8gBltWcmPJJEWkoKRCL2uo+
X+7yp8b6rLLFLJsNlyYzhzQR1TiOt27ybILpYA27kvd0YrfQhV/34is8NRrYvZ/k84k6RY5qYgob
GzsyGuWqFXi4QsSvtzhn9pfFHES/UVCWtsoEKWL/xYOZMb847ZJkm+wJz5KuP6wQQuYWI0Bm16I0
vI3UGQIugdmnH6T+h0jt++Cy9RCwKggoOecC4YwdQ43adebFslvkFfezFcSreIIuzhVr3GiJDH11
1y2HsAWUJ2GmgJEpyX+EepQkv3edXkv51OAmtcBdTWsejWBPgOnTuNH/vWwyxxg8hbh6v0A/ezKo
7/dNWC3XlZJMi8Jeve5CoWMzDZtIPMeTnkdKNN9sOnxqgY+mscUPbUYjKBg8TmPWTubvWM8+Cfd6
5GbIYguWL27brNAgvbv8N7u6AqRm/udRKZqqgho9Jr9Vtf4inyVmfnRQ2hr+nArsk6khbR4gdBzA
wgtyRdMeMiOQUKa1uQae2bYV99RM3NTA81jqZmSpvf5Xe797MBmPJ/qrVZVVTXAQxDu/QqPIrQjc
iHpgTnDb4uy9aNcMmwK7RWEQBjLzAfEqTxMJ+/haZyN4DvpRlX8WnXHRqqPjz79gPkVBDZXeKv+s
/wFICZ21gFju4Tn7sgz2Q7HaYtQi6Px6ztch9wrPQwPxH2QuMviD26c/8wD3fur8g4C/ukBsvYH/
7zNdD6DzuNzUB/EoqMz/tRpxrXOVlAW4w7g29FX56d6QKHVKPDF8AxLgMk8KuW/S+pBDIcddrpri
VxkMgk7MT9aDnJ3ed5Ld7XrovvrbAkvEF2CQmv1ZUE2IoP7ej/X2wyZENnQAc9OaiqH4o9rj16CL
h0tex46Dwsh7j6ZR1d3+6u+GK5dwxq04GTW0rXc/eg4Vu8xWr1qigeUu4+eZxKVTekMgGBKGcc2L
rgXIsKzpDBaSX8noTsIkE6Put09HgwGf5YahhGP+zcKtSXOo4cjfKzx8jtCkM/oNqlDW3bWCY5jk
tiUZ2CzIa+SBr67Xrc+dzbxgF65H4bml32hRvRZR2CZbSAwdQDwSSwuE28OnT0pkPSaOvLJhz/ci
zm5n2R5HXkoagj/SmDUC0xtxvq372gYNPm8AP+ayzSJ+2dEiXTHXmUN1h4N4VhLR+yHxnq3bmls8
ap8W2iiOOrAI/RoMc7u8KhKTdOIX8k6/hp9IaKx90prjmsVvRV6K0IgLj3lpv84GfSoyyRhsHt52
IA22YW+QuWEMZMyBnW7RrBZSBZ/akR3fbja1uzE7uAcqEsW3XKVPo8lDj/B2GOENVu/MKEnJ9R2b
0Cw5Wt2lf+P6YMPqU0X0ef3WaQPlD9B3Edh3BLwcm2uVRcB9WRJQy9xC7GKtcojNJImFqsanFwgt
SLD6954V7uBDdb8QA9Hmvj2kjrZJWDXXHwjbAeJqnGC17CLjE4/1vYbPlPih0rcFQ935lLIqLQ0+
/asHJV5sE3M1UnkvSyjLAZm9hNwSpddRht26GBiOowKjdFav9v5agfZhIfFiTU4Lwtc+xyWpDROB
hk2mTY9mLECCAxyVBiYUjtqqYybPdfVI7r9Gbz8Vhr97PwI+hJOwZcTm/LlDVJpb8JJLDBd6woVo
uaYP87RVBK2tASkIeNiRXojPi+RWnpHxMrcHyLy2/cw5uBWdI+ZjOfiwMEjL/zxKUQb5a0tiRtg4
1dqi0Y/v3NW09V+bZ5y99BsKV9sqydZd/tIeTsNyhI43udU1jfYXbCQMplbVRGyKfifIur6Mk1BX
6Cqxu2vi7e9Jfm+BQsBp4Of9OwIOAe2Mms9fKHonnDgcdppajPjheve0/upW3tXspH8bZYNQZ5S7
OBTtg61HOZ9vbyg8VgphXIxhqvl1Wc4NickHeAXjoJd5hZaJuUuGCOeuVTR4ZVwUN/jRHBzFeM7N
s19f+vvGSE3duhuBYMUwaa1au3FoAd5SixFcqSBqZDf4WNigjCWAqMXh8D/SPf9aUBgbym9OLaBj
vuCbPujXWvEEeWvana/VU/cyuRHVMZGuFL2YlJiwLrQvHzNOsw9UNE2kq/78oU39zUOvtW0QScMs
k86trS/3+bGOk1nhx78xWP4XSGCvNONAOawdplCD7w41SDHsXY2D09t990Fc0QD48X6E4YKEUBge
vyh1uBhtwcRS7OgD8LWUu2YGv0T9EZvQuPunVuxc9ZnsqzWZhWWXhKQtjP/07K/ZMuY0QM8zDqUa
7+d0Bu4QUQzf4CXx0IGdsfKAnsfL+U6zQ3zA5fbCe7pjSiIBzC4emkbhS0o03HN5MVfq6x7zGa3z
upG1EhIHMgdw8lRVi2WJ80DAxQWBOQYHWqvaHSZfy6MiLgn581ohRrasJQGMliFo9rOJOyEvsip2
mmdt3s2mGrVyLeHzVhCJ4qcq8noPI/XLH7EjhUeb34kBW0kcQ0/z2xf/uct8NzFyxZhRz5DJTDlu
O4Dzv6vCPebyFHctiH17uVyNQIVnP92dP83wwKoJ/apSPStFK95Q4b6R73KgFrCiNG9kGCeTGRs/
uFddv9X7hAmN6bYgw2khbbc9kHxAmtXIOHEIYFJKAqV5Q346FoA6ptzSYcz9CSAi6iVs4sgutqxJ
dkmPN8RKRnGAUvBV+zLUyikEaHX2UM5JcPr/VKzrK91vbeLwUvESXsK7tz3Y4xwKm631EL58NTFh
YA73BSwBcLon3kDPoyaOjvL13/FkHTRNanKcaBXUBmtrj51jGfWf7Hy88jqPNS/j/pp37tRWil4U
2+AO73fjRYG3Y25qp1tlKu0VLQNRd1xaIr3HKtu+hIGbrDz6/670wCO5WGSoepgt9IpVPFuaQSGz
/TN7vt+pCDD3gekksBAXfghSDy2n1+gP1AuNsD3ZpZee0xdf330ULUx52C28IdAHnfiRRyZ+vl/7
5s2T/P0tPukHJT1/eLcCXXYBRKmTuvoaUgzCT7ggOxxrflqus5OMnGXHyMsJy+6cDwyVmDmADbYH
i1r50XLL86df9Cew3urZJ2m3Yboc1g9/rbhCx/OrrdMrnJzrAVSF0FsGRpl3CymUxAjqN+A3hwE1
7SRFQGA7hs4YXQ+11f13rfzzFtxFFZbFMnmqWr04w8KVRC5Pnwl2afYs3+KYWGqQ9OjmL03FlBmw
vDO2aYZZFixML42I8Og9nr2MVwkv9oOsmciCpnlMJI75WQ/+Qebz/kpNFaWhtB7aCpgjqqEvKYnD
xpt5hzrSEY1TqCQYjjXw0ccYauKjbDiaVtwt/MLdjak6StLEPF3ADOHJTYtmgBGUsdW2+kexxBNP
ME2PZqYaWea4HRhYSDfmEGF/M/+gZmtsY7PV4wM2uodlBKGYIMN+60/SEOemRmCpsjNP/Y4Yb763
v8XbhHw7J0TkuL3mO7kAjC/3N+hwBfG1zv1WSGlbfq3IjJo+/ZrnsHSb/Jaa5FifGcR4mg6B5C7C
wsswosXKU4QQK9dT7bOmdlThY3m6eTRT3KKoG4RAG/kZtdqCvDVf3uj/p/UhP3ICAmv1SWy7igIv
9UW29kRrj2gL/79RwwoBVdj5CJbeZzS+Oolh/DMOe3I465cDOW5a4eq5ZcAdMN2dM0sGgzjkuaKv
zcYR1kN7ofJKA+pgBtfSe2a7GpCO8w5gKySPDztmgVGrTYrCcm0RsoHP4OqyEwP8yOaJgv764IWc
Hdo25B2IZhdWCvE0kHKq+Z4ueCWJP+W4xEpa0bjceggVIm30jUFZ9tAMSY+6U7N6OWYSsvqYVuXv
2HIkuuCu/VdEjlC2yLNWyyZ6GChBG9YUtKj1nywUnYTMSNiafRpJVhl79WjhTsdCSpsCIZOBRniV
5oAidoYKqmobJ1FKSqp0CBDXUyJDqL0w4JbhQ/5mkDxGg8FQS9zcwc8bH+UUqPAQIi6w0eZcp15Y
l4VB4xJXuGw6n4Rh+rtxqw0GE/MiE6Q8+ytoqp2vzSsbfbcu1h6Sz5iv9C9WxIwMdaYJw20t5Uty
1T620QCnhkevyvJrrHWmJmPDSBZj1QOIohUrjgt1PzQkO2HyfqwqlpBDmLXrELzwACP1Ta176cvI
qS847BT8pf0vfF/Jk2ywr87nK1zZesG1t31jDhVOzUTKwoqw/7DrmbmmplubuWWOm5XeyeI3Y9/d
F0mtVWmWtNwpvDJ29Ze57MTyBSvuyYl6wvm2xkY/BLcMopZC/i8BIv7hloki6lOLZ5uU4D60TE3y
neh1GaZQgX1tvQRVyuBQTxBRzHYrzVSYwLq4ldMhOGoTmB63qVaHIzYDrFgD/zZgtnEcJDpgSraM
Kfv8Q3LCaYhxmYkQAD4kZ4opASpReCdZxzndlrtf3EKQl6dREeHA1PfzcEnr/r6xd4PrY1GG5vFO
ESTvbJ8YnRUpHRVWl0/9BylUL2y8DyBPphjj5aAJigp3F6igl1cvxKLeh0ipaD+HItUDX+l81sM1
qS2sxC9j4SJc098OEMhPzussH/jZ1ddFIMXXgMb/RzX5zVVgTsQeO0YhvMbdKCCmvPaljLDk8b4l
gP5RPMuBKwh89IT9v4xOlDab3LH/EA+iI2LxowfvPkWHbvDZCv6aeydKIYHMwSbj0MNtXKlaF3l9
OzNxg2Pp6B+Qm8DKGJ4Od0kIhU9KTe0IEgJaPWVnjUgRMbiDfyZZmr7TMSmRjPQp6VjLxsaXLEnn
T+MLPt/UfBwyRUd9hd5jxWMgyeQuUmLH5RJFYhfQZMnQCP8bMEvTs7TOuhp4NzUwZCNAhM+UQxWZ
P1MiUwS9vvdZHmANwfJQWUkKeq+SCLy1VYMjCGrAPMax7CoSJgU4X2DT0E30AkmfABOk97DZZkZk
oLun2eZRF58PChlaT+f3Mlsn+5QmRYh1PraWy2YQr3+JlgmiTC9/cb4OTTEAyKT+z6mEnzwEZzgx
IWTsD8wvDAvBUiiOzA85vCwV4h7K4rx9O3V6py1QJykyoTuf5j1Tz/dZ0142rebCCzHbrHWYM5Yh
Q1jyxYsyLe6cS5bZcrCS3jF+05vv6lj/kidJ+z3cpsWI+nyJ9u/6bt+iv8PdZQ+/94DCWe7CKAxF
p8akSoFwM/OQ6Dn7oi9cVmJp0eQpSs05XWzGLypg7/nQtVJwspU5lkl2K1Lo7pTMXEGKeqrEmp6v
TuzplTS7kiT0pNnuLKJk3THQrRlDOF44ds3aAYe/8IUrXiKypFtXHZMlsXBKKMTbWW8+ZkgHKt36
DvLq/xQW8+8wXf0VheW5N3Dwiyg8L0K24cJS7f3GvAJnB8kvm3aMjlt/tmjc3ZKFQDhtExFhrHSV
EUTi4A+k+JU13ZHCFEiVQgJdbSUVlV8a8wVfEeDRL6FR2Q6CA/e72W9or9B5NDabACosVkXCHYHr
khKFWQM2uqjz4FoT/RDdXZaHw0UQ4oRLbkHn116AYaMfTqradDBTs91W5XqNt4Sro3VcQis+p+55
hcyWnism39nsDtFCJTV0I30tTOdrL3UDf4zDMsjg7r+4UiTFk7VfNDgNbERCb78oBSKShvgTz2WR
kedJbMPo2As8SNV8pU0abqNytgRdPkEb0bGOJQ7yKftUIdcInrhpx8ulBb4gi3K/riwqwhFODwOp
s2emsNQatyv/KxoBg1newMyRk9FQTvbJO3FrMxTPfGoRaW9HAA504HIATfopOHF5oYhZeRWmze6J
nwNuLNAd3dKtBlKtFawAyf4iG0sI1o4Sqxrgfc4Ivcc5DtRz6reYxanyCPvqyot7Sc0Qx+/L+qQE
/LweLE/Bcyo4Quc5MophLBU0FgRmbPa2yyp470OrgWpGQ1sfhSJQkl82mzoC8Xa9LTTSX9djQrE7
B2mHpUJ0u9njyTPfdD6P0j/VGgBlKh7A1TGs5u+/yo8iIbpgXgLLKyavJCAYYE8Llqb6Di6h+cBm
FmSBmhJnV4Fs+k1hWthOJyeml449AP+QH1bRTNHSuav/aCn6++tvst41rTs8yQwfSxk4IoHk248B
8rr1xstSRZBNGba4yTq1Sc4HRgKk/UdHp4B2yBcfvedI6Bw3LZ9UVPFtRq+Zh0oUmzcWoKZw1812
RnrWsUnX3XVVq9iRny9rsv1nTQIUtALzEO5IyN/0gPnUn4q12O5ipDsMK1zrYXQjiQGwjEdWFgu1
lTF7mDAEPbTn3ODXbrMiK3SoTYr12ME7JgGh3NBAY4NosnyI3OF04CZUMUdbavTVxs13JeEKI2fe
VNKKSTDKUBIy002Y5rozdSS7+p05QS+0oJ2JTaqWdB9ObWXUuVONJbI1BOfSgHFk0zVQ2kGg5kH2
O/BLrrFbxeJkvwszmTwGgeg5kRJNdTnwx9z4mk0sPLALjp80i4fV6kyWaQ/jpwu4R5I8JuMd5ASF
rBkFwBI71tJfNO7W7Ap/zTXdhKlx0/tTAwcPPcY7KgzGLyOE3BIeKFdno0WGTbwZ0jlAyTwZCvvj
XDcythNIOtVtxajZHIjDiCOcENtFjZ7AY/Uv17d0iEQCF2dQtozCYW4D4RWnb3ofRM/frtRtrxrS
3K9VU8LHEYST6EomB8E9yWD+JGJIWwMnanPs5axopWo0KLf+Y44388872T9XnP8IHX2M1O3PpbsI
5rezDpKobqlqm8Y1De1AcCOSxm9S5aEK7lpi1rakQrX/nN2197S7OHFsJJ2WGssBuiolqrxocGna
TdvpD/scvjCK9AFe8pHXmRAz0bJrEaD3GavJnet75S5sohd5g+vhVcAxWztgdHXpnFZn1ZNR9UlI
kARZ0QzJME91K1f5cflKp8SpZONzhSBcsU/OidOxJffhc3ZmSADNgoVroamctsmwKseJQJXdnXgA
3/ofBV/I/vSopsuDKfVA0VTp+FxizOjK7CPdu20yg5SG19j43+nGSAvCvj+Pry7VRqj+4HeAKnuK
qcmuPxH/hiIqgEuGkMUab7DWubo3whqGsjzZcaqnTL8I5g2+p/SFX0fbVBK2DoWp5kridX/BwOmt
/NtmM2LrLx+3RucV5LPEq6+SjlOg6WvkFXbXBgy/tWEJ8EWsJAc/navjGsmy2DARSnT4YfHf9psD
RGutyuxJkjpPNY6tWNkJLOJDBDIVZnZA19M/EHhy5h8LHgAgWWEN58yMlYLC72PRdpk5Y8D48T8f
5ff3nou3s194n6aBt0+oXRbeeJYmCeqNYGJRDXmZK71l8sHq6BhCvE9WTznxIbc+CupTS1W/ySzv
Gdvum439p92x8TlI0Q3kIX81CkU3uDrj/n3yOnHkYpwClqy6IVJ76Z97dTw3NKCj99AXHEhXMF9R
p1FAl31tIs/49KS6MfiHKDGGwAsvIu3RDCtD3nwJm2wJTqiS5DzEKaitiYFhkyftU/DRTb7WphJQ
ZArW9mGzLlc0HBqOkW3nJCIpU9JL/sIE01vrSvAf8JAj7FtGUL3rV/c33JdVuGAwh1N3hITFIc/8
s3BnkRQVh/s28IGD6bKldCOgfpvPtxWIpowMZlc5rqZYUf6f+c26DydXoMwxHdZ2g30TZnNceohR
PvCtFBi/5fIsh2dQzHOgaye51EiE9gp2XyYpdWPzgTTQvNM76sFLOmGpD66eZypFHfh4b54zgais
5uwmEx6+c6PBaGAqdC6cn/w595nhghxIJWeEd82+BSpcJWXTIs19Ht6/8sRd604xuxBbsCRb74Pb
E8S96d9/7H7omthmufMaDUPrACnMQcZ8l6IGMaeQe7oURIVCSxvjNC3eMBzYzJm640VRyl42uBAU
TdGWuBDGE5iIrpRf4AX9z7NEB+UlxYlF0GZ0o76Mc0il0QBXVQoo+bOLi160Hg9vs0+PFZuuDrJQ
lQ3aQpA7Ifj0W7GG+qvPZgW1nV5prmaK9qGfgWssWUlE4nO5PmsxkMVWUZqg3FwCEM+Rj+ouhXLC
ImdzWYMhsW/kFnbiG2cvdL92wPosk0sczAOBTFM94yJmB09c0v+CMHcfVkkrqtbFkCA0sN9Hx90q
j4A5jc5WE58UdX1de0DmncPnuqxJROnrAo7E9k42rrl+j8p0TYV2Qud9qerBWBlY/YKK71Uz/4kk
/U20gVSxY+pLNi5u5ENToN2Ys3VCR/WzjjJM1fjmwJAi1exdZfsHPvSznWX345g3aPp03L2/HKu6
vqn+2WJ9+l3YF0hBPXho+YsUZRAyt9SI436jbzoUlQL29qEiyIxI/aUKPSroNH1vovO3cODoEgp5
P4+5LA3hj5OsPvz/Z2OmPjswOBfUYKSjkdJBb2TSwppjNIAxAdr3rrDtTpAdP+G/6o6AL8vMr47y
Vy6KKHlAKjRqFuvQ4bwbOs76YvjPbdSUlC3CW9fMrCGBnaIOPuyzEpoDEPJODXv0UXQg1vLJrbbM
BkHCoFJ1HSAqYNBuaUt7vUth64z+JVBdd23LtZDe1Yfg7wiZGcwL8ieqzcCw0/KHZ5FCQaFmzSVo
Tm4j/LA8QRvPj3ps0xpDVyOENwEWGBX1emmkvMWC54Pfnr+xkVra8snYX+fhpXynJ9w7RZGfvxUC
yIN8ymHO98NOpgAvZYW1qmoXn7khBnhb3TperaTsxnfOMJRxvYrCVfPe+MorVCiXrc3d6pdH+3gC
L5IZjUzHF1i71vWylLOzUaEgw+nw/uz+WffvRA/AV3MtSgoCv3sY5etsdPjIEsx+C8oYTvt/DhZ3
mnaqnRRC87B25HKU0W0ExcjCA6NuHZDE4aksLAam66rPsRnbKylBFHWnVeeDgfLTRzm8Id1GRzwG
oUWhN9Qv5OioP27WfuBhLjOI3Ut9m6vR9M9pg0or9A9JO7Nw3szdozaWPXb7iDq+1SXjq6R0w33K
vi3WOTpJ78XBKi2bHfWYi0rbXhV3Wj8SHSq9QWEQWgiZSiKiIPbLnJBRV4NTenUY4wf5RqYB7EcI
04PLA3EpWJVyIKGEYwwdDqWCw6xbJtVAKc2jb4YRWfm1OunYSdRZoE5Dh2xXlMyTT2KRt71l98JE
hUiHtZlxNVUQUi8eVxq34IeQarSyL3PwpuqhSBFiUpsdHdt6D1pPUKFhU58Q3NRjsWFdykOiecZj
4hNPndH5oqpeMgrceJVC3Wft4MBuH8bu1wx+496vyQRT+W5agMYnH9ZRxSqliNrgJy/caIw38vne
PHWjagVB2VFhzAFakDxW10zsLKpsaYzxa3jSNu5qBl2eJxkaYVsguqOTxmBiXeRThM3Y/tFjmgEE
wYGW1qCSoaFc5DMb/t3W8GxP8gTT1kSzrGjQBerTfKCLa6GumUYLR1Okll1G864Ej966jBE7p/QK
YdDC0By4/FAa/RSEFbQShcVNeSpi01TpC9bDe1p1PFyHDLMS6tZfhPvq3l5pPa2xHNc2ADEjVMDD
JSrBjV7oymdSHAqaDzvguPu1z1JdfvXMwKpEogaFCKV0qDDz6yro6Lk5azYyVDWLq9jXcIregdyT
1LRTQkBOsaURhQDsZgpmML28zEmYXx8fwoJV2KScRob58u3yOUqZx3ctFRKCrwDUQAazx+ZH517R
jKyDaAeWrNV1QBhp3CXEgDZaUNbjR+SX9hU/RGQVdAIzcxGoJcE3WDB2Od4TXrTfS+b69SP0pZlG
stBvX+p7h+HFbNMMxNcyqh+AV1qocKjQFNINnZgXR8ySciDOXwmVXNECHeZS/9VjZeTdw8tN01w5
IQhRo35L8E1tc9NziQCGcUeDzgY7IE2tjktfCLoYRBHNTYZmo2wAi9ZUjG4wE11FVQyZrklNs2fL
ZDd0BBudO1iFUArMNv7mbGsqDt48WRP8qC8weqpkPvWqor+TILGHx9+tD/GmKpgS+szTEzNcvDvL
gxqU8KAEgvYWTjkBImZNcqWm6jYSbrkbmQsik5y8Ya8fdGwChgDepvNuwYfmZi4Hx8xqx37864Yv
lCE/QJk7/O87mD03GuZ+T03G+3LVpNvvCZKZmC5zM7CvD6bsJxdXXwoKt3tKodM0gb76asHDhlS1
HajHGNKiCzoOCj9QAdrWU7W+sSJqNkGh9x6orpwlrojb9MQeT0K7rXgwtaKynEWbiOoyI1eFsM1t
iHVHsiXww2UWV2wde+bRafnTNa0yBjdMxblNU5G+PTVJFSnJuaNinbqlTQKz1MIxMKVffnNfNyiP
wwfCNY5X3NobjicqeLqHTlRR3a/G6HTZhfZzWenrDMupTXclUJVFk8989OW7TDEYypj59YL8GWnx
v3rno6t99CfdXv4Bhoj1ft3Tbss0axDp8/F0DsVeJjArfx9YmOexiZ1c0ferq1VeZGWZuVOht+JR
kALnaknxon4Li7XRv6dLKe9FkZwAwaIodrpG9yvZoPQJ34Gby5GvkEbAZ0SoR9Bkn4+muK7V6Qwg
5TcDWScvLMWYDGQIjkKyEW5AYaMZ0MV5aouzDTSs5fMsy5fUvlRQUi3gzB7Zvejy6nr69sSbea95
yGRR/Prod/COH15nRO3t0E7t3tNmrjL4nV2Gh5nS22SPFIdYKb8DD7WKCh/QpVEOJWtwd4gd33tV
JjMUuZdgSRkBZeRE1xri09CwqCFHBckqpxOr10IaLNcm4OW4uF7jSK8iQ/D7/qP0W51sDPkuNEW2
GYu+RtOcyXeVKw6nX1JocwgoJZimEYGFnr+8GSmt67b1K8vNzNqaCpL3DTs7mG8hpoIUPpEVNmG8
kaWfCaqZR8VscqFqlyOFecM5JaOvpcyl5G1WNI38g7Knuv0/KzvZfZT0C5CSc7tafupViOTtCReJ
8VP2ceTF9ZF5a2v+zhxpl5oobL5or/sjSiYpPCYp7d44nR8Wzrwq0+jHccKFgLLuh8zXSQmOLX4Q
cWHrm/k5ctGBgoI/h/UfMMUhzBKrlRnNTGB5h5f88/qQ3T0VJNAuP/Q2aHGRsg/r+/kcul77KQDw
i52QUZwyrVqBYA4NfUoJ/fiQLuZzPEhCYCiiA+OhCvP89tL20++iISHIlBXc5nWGALQOHsT+YnOi
U9MYLjQP0wUEz/4MZa2KMmIWkWwpweqyB273Q6EHzLMjFW8cWzWw9/2ezgIWU0Ug5E4G38HiZBVF
EUZN/2BwKjTglRJDGG/fJ3EHQHcwAGfov6SHBry3xyB8yK6fwwqU2y8Zh6TOto0rlngIEyDRYYrb
9jL0shWhZ0rXfFPJiDZPRcWrCp3ugrrbdj8jj2Dyh2NZUFqWtikNGOykqIOvwy6LxkNPDO1IBIOU
WqcNEscG5Orkeds8EY0ao3Ti5jAlzXlTBDPQtS95/23kIY4KbZGn5WpdgNNTBflKh2zXxwVKr54D
TZGiP/VxsascQUcAD/JJpHWyWf1umXygjYdHvSXCFZN5j+l4Euz31NsCZzw37o9d0u229Qya0IUi
wiLj8+0UES4h0qwWDdvAJ3Ik1osLMfpiM+nqIOuKo0C12FLhcd9G7FxU8BUVBLb91uxlL0m8STde
7MtruDbEXMhCY69iYvlu1ScUePUY6Xb7aquWMTJ5afXRH9JOX295x0As4zH9yreDmvIMWxJB0T0n
hQWPFu8kBWEwLHdijRlSRjA1/YYOBYPhr8WSnaVLQOjv8y1GYw3/p+0IUqTzW72vqqUbM3oNUM7s
49wa78GA4et7na8d19jFBFRYpCiDTRo+Watt15rpluLDizBJtJHMqjKbeXlNLKgmncHFo8lWSU+r
WUPo5mw+afwmQ7uAGLm9VKKgYDFm566BBww3m4Wy0I+JmVz3zTwVyqzVhuCETVBY7aAylQ3EZioC
TrrlhVMoUsF69pEh4QQ97EFlW8F6zrjMB+3knbgBlBs1u6LUnVyFc/vO0soEUs1dmZiIvc/3nRGr
+XZ7414mQn3OCu3dA9yVAq+bkpDeOBUy9RkTsTlwavCLfCcI8grptTp9LDBb823+3fBucmoE+TYx
60WTDwUcvm3Z6ake2pdgf+muIDT70AamlFVRSrwgWbP+jgnI+WoI1JIx/wHn1ciojNT6AgRhefg4
dlqVeSOodqorJgfzYzzgc6FsHipf0MS4pUgjhGHNvDveKALW3bir81TV9YveI7m7AILxuRF3SlUy
6G2wUPwmJ+9ItWu289x3+K+7B+jeEg92oNXgMNiHlPcTQRIkXaQJ/4cJxPVElq25yQ0ebVMbRLie
Gks0akmISqZ1wzS867gPZU1Pso7J19Pg/wcFxtehPFxkOGOL+BoSlh/g/bCKbP0Dipj4GW4ljQ2T
KWr7B22EdU8JZWfeJOh4+adxQ0P7QdZ4GVPAjxe2xrDrH/hcqNGx3wIHwtxRhmKbCFs6c5FfT9Pk
u7O91oOTJy47EMsweDoTKdePSfTdgVMcD7omiaWknCYs7ugkgH+AZ+EFw/GzEqPYXuZUc3sMQUJ3
B4qCNCKWCkQDBzb/kj5ZzbGM+GTqw1w4b6p/Jzsm3Lx/Z5Cst9G2Tmw7TzwCbNeW+0RbFALT/RxW
2fCl1luYMHvxH6Lrl4Er7ZslOveTfCQMtyib0zPf3BP8deObEtfk78d8YYFK3kG8qXQdl/RB5uu9
fx0QP5qNtMSwaqmnvU7qRHQq194QzYytZTONrLf8uu0JEBANor45TqSqR0PICBoRjl7i1dCb7z+0
iLjC/wWSvakVjtHiIMySZyxKvPwBbi1buYzOssaRrzFrnVoDmLPTE5pS+4YgQniomSKD68Kkr5X1
7QFLPI5Zc55FzhpWYfX80dOwfYRhwYlqyWWBdHrZPWuHksFafJHVdyoMFSMTJKfY32yD9X4uXyV0
7R8/eKLhJhkPxT1Qj3ceuVigOeZSftLSDhZR4lOjgiGmn3IGy3BblnBMTbzsiwqa3eHJ0eEYZZqD
nlDcXuA+TtH5LIeiuDo7305lXmUpvjnqfI3B/y7zrkJTNA3gALBF7zlBWIkRuxn/rePukel7VTmq
vRNNbQb/T9tMR7cfGq5/cn19YSaIdqUOYYZKZhIVnxqVlSIL+xNBe2X8LKDFUDahGC99rtJsY6Hu
KP8cQfDHBIun2v/3n/nzrAG7yNlxfwZEns0tiwn2gi6sN4q4PSCm0V16Gb/SiALxqxSN6LpL5siE
g6w0/Eo5ojKh4x4oEYR/PCUodcj0Mr0DoQc+dw5k7/zBVoFoifDKEXGHeRibmpJB+8DrFLdVY2c6
nMIm0y8c0LI4apANxpKPPDQD1+c5ooozjRjaRDO4StCYPfFXB+mq6wQ31zYBY0OPDtjmjCM7dTi9
/890urWOhKOL/zO5rXfMblgDnxuuM1XX1moU7lxvdpVP9AsB2jspnFPs2MBY5+VI0AwgdbD6F3tH
v1L9fdrdtNh6u+CFPjCncIJIIaTlNw==
`protect end_protected
