-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XzKe2TBjr1qOPwLkGCzyaCkWf+jA3txY2JzxoZqpWLrZcFxVov2mwaJAyGxgFUkHImb6R1jqnrRg
Y7zJ9J6XbU3849gh6jhNzvGM3HbZW3lnKE+L7pekYMgwhpUDSW8wlRTtWic/gc1JKFSP5c+J6Blf
zxktc2S1l11RlqqUq1B6LNiK4CI1/5418Ui3xtE+0uPj0fQ6aP77fTAuWh5rCwfBkJX2yFVl6P3R
/5tCZFLu92zsgUWTuXqy+4SXf4fS+Eaw9Rv732497RGMvnEsXTX5l5FVN7sIDcxW7LvuLyzC/K4y
+pB3AxzX49MTiydQZOoCU6ylED6hAEcOnnzFLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
w+0CAM05qSvbOCf1DmqZ8k1/691wH4FYdZTryiCMJVB7nyJfbvBbEvdygPoXQ4RFKSzyUPKb5k9m
NJgXd4RV1lqOiiomnNONRzZqldNer9ZIeWC7mmzvRDMHd/HQAYLroPcQs31XHhw4Xb2UCMQrj0VU
b6U5+OLfAg5OG8sH/SAmHSHYMgiC/SzYm2aSFEOPXppwDJMDYMKlUVydOZvvs+e3lewsnIWKz2qR
y0QlXM/cgM7AcmdM8JPm7WRw1gvHhiiziVjXMx1rEgzrW6VY5asJSPzwsr33SSvucACC1gmDRPiH
fkRpLaDNaF7xe2QqbKoYu5Tr49idYnrAWXMPnAXJonsIrz+bouacGuqc2F1HHfdYz56qAGrX+HDz
u6VHbYLotFzeqG0MDuCW+s5dm7R6ESgrlmP9P3wWn5LUeXzGw1vK1hO4e/r56+2NvDlekXn/MMLH
JkB+9alhlfl8i03EKHfUzjtBUIOMe9qD4eDyF2WC7c1Ts0yeXDwAIRjIm3Rv+KsHjsQVLoIdsZT1
8jyCLiBxp6vLt/ou1H5Y/CNCnQh4U+jwii+2FWv8ptzcDpl2tFjEgw/hiD6t4ON3hhikGBwUarFb
MILpL+vBZjYkiTcrBo6axOO/TRaXNjhzKjTQFHxkSUx3N+G1/B+qPD8edglFG27itBhduSOFpl7I
2vjotRAOGSJ6Qf3lbbBxqIj8WxH1/zf6kyyF41NLmk579dOkA+nQLi3wtoaTY9rNvXT30emsMhL6
N5xRsEmOhriTF/KNtsXMbpmkd4Vgp/5xur+i3WooEOoLtUUtm4iyUQL0T2fhBNqHeJEo/EOP/wS6
17OKkG1mbCpciqmIEKzE9Kgv5mpSy401JE8i0xJPIAUEnaNbKApMRzBmgJ8Hh+/iGYpeM7shvxm+
tYKZgEALPb1raMcesHCLJMhGEomF0LgByFhm68vGcQN2T6mv7gTWUgatYAeb6vJZg0taiuUcL3+6
r7AB9yxC3gNK0LBd1aUb1cJUW9uv76AQn9EU3mEwyW+3GggtExduxWYWeURnZa6ZZHGUO64MmPRA
N4TmwamNyqKotVwSZhy9lyc+TRhPRuUWUFvkSikIm4ttn7Aozt/97yMhf2CeA3MUsI458f9dPuar
BIoDy4eu0iD1SW7ntG7GhxJNJpnGGglFIYJxVruiAN4KlQrwyS1IfRmKsZWYhGjn7JsO4D7aOyjZ
uP7JcVnAmLW4xOa+wcfx9NtH3pAJzoMW7qg6KF4//40P5boeJZf1oaLYCoWBk89BuqitE2ncuIvR
SYhHd9YlQzTsjnFZHbHePLB44Rjhu3J195HW4ZunghSD8tLuz8z2hL9JfP1eWKNyumzSG8G4fnhq
tI/OTX+1xYeaBWJR6R9ZXrJo/wBf/4TJpgI0KT/YisptRGhTAIh19FcqCDCQg8r0wE1tyuQKiv7C
wJb0LpODtOzgNVwFvxNQ1hOcVs/EApbf2CV/oud/cBJJjo2dSPARUsFR3VsM/HUq+9C1F27BTIUs
QqINO7Tpgu4ygchVO6SjlgH0om3bd0xJ76IrCOTcY3LoquUXFsJDbblQih/N+TExYw3qPvwjUCSZ
lXtKt9p/yS4JrenlmPZO5h2n45fzcHTuBFEY1ZBDH2fvkusavUw7hkol9fZKNs5I3bV6+6bYPXVc
HVQyNUIet4z91N2NYicG7jB2LhvvkRqnOoH80zP1HYPdmV5yV1EHGci1usetBwgMwkS8ZDa005kd
OfbivFZAEy9jGNIQO2nRn0P/pjMf0iwasxDCsCtXmjoboB8sN9bOnIQnj4Lb0iz6N/BSyMYtO6BD
dEHU8AzvSQ9JO8lnfcQJAHDXq0MjSXw8qh+IqHje2xWGPxauLCZ7Z9I9i3GSEHU6/jTkDvsm2GaS
TMxPQNAT2D8d9+fsa/2nKjxFHpg4/fawXH2hXJxJUFxenig+atNzB2R8KNIScrtpuF3aqvddpeVG
ik4XLmN4JeJrGiTUdF8TdwcKQEqNGV8s2Aab1g0IE3zPtsNFpRXzR8m1NHwkocsovt2/GpzNi8c3
j0uRqO9kqL97gXPCxEkl7bN1p/9GsK+bZUMa559cY4eVT47C9sAAQGsbDtspLios5HiOrVb4YnW9
/NgGGs2MBm33i9i+3fAAS1z5pAwHFDr+bfgv8j6X2CUQbD9EwRYcDyKIepBv7KBkuKOJoxiGYdd3
bZzWDE4Cpfj7z4MIknA43UYAFkTN/aAAtL0U8P64KNK+M5b2reY/V4wHU3hn0hKZJP8PkVRP/4iP
cRbXPCBd18Fu1AM4hvIsnB+nYZxfuvJ+oAuIj7DxsoJDop307uFeEe6rTf/VFN9fwPjudiGj73Qz
BGTlAquuLaGtytpGkM+iS+ECHY+cfnXdG4prfDjCC3Hv/RvLqeMJ1Wba5kEqckqV0v3zJtVAyzV9
JfwRkCIaTLnMc8Crdd5APgdDETrKduzb0EFXKLdbP7mDidWrTrGEe0WdmPBuAp5K+MPv028gco6L
pPICaFZDxH3lGF/4HZUEJZT6TSX4jMGdrWcZx1nAX5hbYbh7bRGd4HjsvbB3fy4nTIQ6bluGs5Ed
m/yfQL+pYzITtLxMoSoujMRlZVgXDTd9/nYKDDKsGYd4cIr4HjqHXPB+lSkEkN/zO3jK/f2Xx8cd
PQXS52+Afp/lAVUfYMXttPo1065JdPuIC25rIQRbnqEqukWF/9qBkAnzzVCgiN+XDegTJNnSTTwN
mZhCLRqMBljCf7HmG+JswZUB40lRrBIItWxKYcrJ4QKqQhUQ9ujpPmkfHgpCAGKnJtn8RxFMAX2Q
26gyEJ98I1qbuyP7o/HKm5yxjCFkG4B6Q/OYAkdSn9z1uAY0/ySoU9YiRx/+Xk1DSGHi5pmarNuW
zfy30CDOYQ0z9I07S/xG114T4m+IbJLUKafbMj7MxkM190DB68UZNZL/+3OlW60ZfHMXgWZhh/ot
fCTy0yXr+n5TXrtQAnauEnCHprryAyALX602C4jTXM6ClwByjgRRc+gg1XwKIQmg31lyxVuaMXoN
DWMLaOJs0BZ4D4klTyP0yYqZ6CIwJLXcGAV5WUPkPkqDN7oe+/P0WEKwESOUrC39YAWT/1rHcQh4
G0Q+ftN/BN1ytwRLstf7/cfP2u8Oz0qmUMyI34HLN6bh2HCvLyHfmpk8itBlK4NmA9qdkbbMfQKX
+Py5mctxe6DbSlqjw5uobvmmrARi1xncIwkOGddNpPrp+6YJyon6VZhn3qJ2POPVkyQr9Y6oSd4J
QniGtBFOSjypCILa2YanW7LElMPU5Z22nSenWEqz19ICaq9/UypfbtP+ffP3h9fWY7ObCsI11sgL
QDpgBd3t19wg89R9XpM2JUJfFzPpC7ixuTkIppl662qH7284kU5uDFtkPGHnSPqnStLge3f/9NG1
/2BUVA1S2VUkoweizqR/No0pEBdHFT1YOS0OHppta3X78jVdB7ielFidfxZn7MNlBxRETolVEH5j
9RZzTu3CKnJ4IlpEe47CwiMluVcM1wN9pEss9FFVK4resEaVXQZ6Z//ntzwDMfOlSeR0+wvsVUrr
f8qLvqnd4TmC/45YcM9c8fK8p9DyCeQVq/q3SySf5uMgSXtAMLVaSZOWU9QTYet2oG7XXfxJuoqD
a22v2Ab5O+by5xcMrRo7kukUkAwm8h6GnAKVEXrFtmSP+BTuWld34LI8b5e5SYBa0qFUvAsC7wJj
94yVqQmBHo7vem3opjpigHez0v0EJg18g04WdBg7Q8f5Ns6kWVct8UTRJOK2sl2SITYRQwPS16hD
z8McWetujycUulW6jj6G4LdSub8imG+z3RXx9uMzsSuyl5Okyij43E/ZuGkW/+/Ttdao8NdWKLfZ
MMZZbVqAGDtnL3dQ1D8i16NiMk+btXkqqx3jZ6GtxeOMjyNhhCUz/PAMt8eed4orhBV65whHT3JC
i/+2+4MLs00LATpm1vBYLl/jDvkZIv24g+LNHmiGCK/6oUEfvX6TsDckwXAKi8hko2NVZ1vGP+h2
wlx+ZF0MykcjdRwgWnzmAgE4QIdH9w6q0ebzT+r/ir7sCMlBq6PIC6gE1jxmqqoPjljKt67VMXCS
0G+MtK/i5XkeI+S2vShkNyvcb64EtFbWoWqfmZ1VEO6VyL3DhuT0Uv6zAwmQOwL3QrWIhBF2OOzU
dDtbw+c7JlSMac7p5m6TnQV1b7GfNFEr1He+eTVzJlUFXxhBWZ5/qintY0dMAUEujmq3BwCLTceD
jrBlSjunrHTFd4igWyf+tGHZ4H0KIfbTrIoTOeFrYuU6xAA7hhct9vVI6oYnbJj0WZfyZNfJZ4ky
+ARs9NE1Lp9ewRbz0WlnN0QSzsv1pGQkur26mCJpGBcVUdxMeZ7nOQKRrRZBpwFzxj2DE4FXn+yY
HcnGJTgtJzgR8ZkWhEPn6Y27+AKOOWSLalYrJ7y3MNrE5BY99QqEjbmvX1/5XLtoJjkk0jq1r0RS
H0rvQ/ojMTqr2WmdEYJfVnwY+4/bOCQbmm0CKo3mG7GlS3YRY3VN7Ll2yFYWDrWpgVkbOp+J4e8T
oKgECcgHxZUks6FAb0wH74cWqVaLfcCYv4w+zYno7/L9yDWT2Grdu2B+OuiiMnovU3NlGUlIE+vX
gMHFGzYI6LxcKNy4DRUXZHWdI4Xzf0ERviQbc+5Ye8FvLf0YVgyJEqmyRDXbscWFdHb9ZUWOkPBJ
H3ce9IhH1AQ4KwAvwbecZ8AfTDTv7mY4GDxhDx1JaxJn6yniTIeSwWYS5TeTsLU1yLM+xBvzvaUM
sfXsxdq1+VqPZiO5MWn7iZxppoTvpgzb/bDQPdKj5Bpo4ffJiKrxMuSYSphkFUI/i0RNRa7qTLu8
szjtNmcOZvxUQCIJXmA2EtkeFztPws4STlZH135wi8YWjpLuLBqRRaiNNgx2EJx1TEy4wSu76pDB
k4WVXvkbf5gwSTCyuL0jd9AWQUe8X/6TyuCWE/97uNugQ7YJvRsVYJbk0dnxeV7OeLkPeFkVv8rb
4h8UO1H+9hnNNJotebnr6QhcEYwfLR47gIylWXJFHUBcfqgORWBBRdDF/C1et9/+rIVviX008H8w
2OydWxz+6/Wp3l3mM406BiPSx13MQ6s+GS3AFaa+qr6nNM2C6ucRBdUieXmgsN+rpoeQxpGYU5Q3
BjfjDcAZKGFhEZ0wzDecI6LxZfFf3kMt0RuEEh6MVKfRfIC6dObKWvTgj+uPZs/Fm1CdKyOd2jVL
YWsgrm8IjSmwb73T6sJnj2oGSnp8WE+j3FZL8lfEkb2n+i4U0jUVQ1DirdZquNXqpTL2roaSvAS9
INvuiwAwxAPpT8lk3yvJ4rwvSy1zlA+R6YA8keQAjdwON4xFk98q9TyYzUaGqBZEOhhvVX05zXDJ
rBGFLUzAXFkgsVW5NkoOFPxanLad0O/LgelNQjWbxWbQn7OshCd+z3FaSAKFkTO8nZA+E//f7X2v
ITUIPibltX30mjzdfksxlPLrQouGVqQcqZQaJkd5aT/Lf12Po0TQlLNZ5VhnPR+6gHJjlsSD69nP
dz/vjzV+O9bhD6z78sL9Di7+L3ozHQWPUT1yEL7v1hdasx1q5Ll7cRZRcV/QuANvO6qW3Ch58hZE
Si3BGhBkePR4g6x45etV9To/zsmT0Tt34Qwy1BLmpWGgips4Kd076IUQix9sCpDnEuIGp6iDJDgJ
xvLiOai6Eu8GNA125S37kGdu6N6Rpu2VXcizva+NFS0yk74TjPMk502Db6leoTotjBcw1GHDjU4f
9eFLZtU4g6xQSXDiFTujwYHy6ZMqWfx7zUYndzvaY0ydbW9aCqwezwkP7oyL7lRYnTVJRNOqZRaQ
T1/fYSrfFpw5pMvtq7pezc6nsdANLa5xRmL7hjj6Tlke5DZuvBtVSFMmhh1V4M1Huu74bLSi8qYi
OrNlia3yr2yN2wfmFR5J0LSVaJyXQRPn12yPgQaLatE1/Ze5MoJboVL2NS+st/IFn+eKsNlUdNDt
UzE34fgzrwv1eSfH5R5cQrmTHQDw27SbxlqZL5cVyp+Ucrjc+8cVsac30TtxX4sBqI4NQBygf7Zz
nzHsk1PzImV98TmlZk4/+b8bSSrlZ0q1twS/yZqf75j0knfRrtsoZ2mWL7zVhimIzN2lW/6DOHdV
UJ+X9WU/E7odCGrS5ay8xhmTmocfCdLxPALEyQBkyrjfJLf9tqfyRJbvMM7UZtGNTNRFTXhiBGEe
171TmQgI0OFhBqgthaXF2f2DCeNjI3ZGceSZ+/LOurudLwTwzelXLXEnGoJqupvxX/ipPk8/0C1F
5/C233Lpe8yT9x2813fWx0eCDrulQ0GS+5Bqu+IKVTT/uy0xyFMUsZKCxEAUm/eOtRfZ8jTr/2Ns
IBpglISBxodP0ansSWSjlMOPMAypt+E+S93iZylGwxZrp1lLGTFDYGIqQFAWZKHLRNgZCfLQVCLA
xxZQBX1Who6R3LVg3rKBA477cDCaygKUJ+ifdQwwFRmjkZ9QeB5qs5s63VbC9PO/1cxDzQGV0HzG
LQX03AZcfCq8jPYZW1M2TzWQFTZfnEySZMyddNa8lvE3v5FdrTWLMGiZZeLE+2lhmKWkXgP1exHp
nDN31d5s8asn8CwuLTiKpLSP75zFYhLwT2MBWm8cqWhVj522AvuBolIBpDUY5A3qnFjPTvgyVM7k
D8OUiiHS0oBMfpUJ54FsQGeBSB8aVp4aIiIWfesm1cgq7otB+XPeA5IsXdSzlujExkPXkETl3Imc
S03UvxSLqf/UmGzRtJcWphd8NampfiaOe/l4gLqZCVZvkFhRoRUNuRXoT7bfl1y/enJeK1hr21TU
lia72q3mIhS7Kxg87aNRfxOCJIMUXbvmkzRJzL3Gt9v6zXns5cAeocaloHSweL4pGZbkejmXMyLJ
IFBk6nBU311+l5J5xg/c13uhcFaORpwWDCUCWOXiH/ur1N43z1e6ZYEZoeW3em+rPcG5lB2tIwbP
DwEI0m9DjrRUSHXaoykx0ycLAlySgItsLke2sjg/NwlpYOLPGz06wjM7uX1jLTq3mZgvq1u/wKkT
ZY7cVMet4NFM8PhkTqGSBzEq1L8xqMlrPbyhXxHI7qy3LwwxdJ+IgO+9xdIl4LtDY3BDwhdb6HeP
zjly5C3wEUkZtk7YDxdyANt1AlmnnMRV+XkFwRskM4CeO7R3QeB+dQAjKU+V64/EVfivv5KClePu
SDvy4hMC1tlkLGe8ic7HR/bfxc4yw5PkhkNVgQSUF0sQ9FZFo30WKpUEIga0R5KkfxuA5NvYNxfr
+jVQwj8DCEPVTkdM/SyIz+gJtAPOhsSYcWWxMqnKHPxdJFQqN+L7wgWxKpW1GboZ0uZ2lplN4Zx8
QotalNZpMCeXqg8vhdv09d8myq4Wp1DwAuzOcC8yaghxvpKyl1Fe67gMJvvE7t9Tkl13QlVDNRRQ
Ee6RRcEaTEdp1v4ma3B/epBTT6EEl9EbgNLj5ok0ZUCyQtYQDhfXCPRKSpCGS1nxdTpLC/hz04LG
tQIWmOBUd1Cjf3H3jYXtF+bPHx7AcnprBTM39lfEJkPudLfPpxBSn9d7fUtaZ4cyzHtWuNoee9rL
4Arz1a8c2L2z0xdAcY114EO0VvkkXceSC/qNH29myEihvAiN5y6D9vBMOdp4yNzb6FW7YRaTd2SC
RRo8NpoXMe+X+faDX3XMx3qd/zXBPXdUpMK1bBMrjj3fpDuT2RT+gJh1efXM7lneGnJZfR1GD+Xl
+2F4IXtyCFMpZx8tXIUQ+jE4oi5Ma43NxSBqBgZeJeT2tEG8fT53olIB+d2fmEhdFRSCIAgTJtfT
9v4QibwE9SVU8S74htTWYKstChU3cLi9qluG8C0indIM7Q4a89MJrfrw1LuDblu5+5tpt0Qwp7UV
RjZEOQkr93LkpYHGueC9EpA7q+9Z4t1F+1s58kkciRiyFFY6OdVn78CS1yQgawNTSw7yk0GTqBYK
lfRFMSLkhx+ZjTXkTrGTzGT91GlqaXGvOCdBdnC164mfixdF7Zxn6tIMq2vhAj0lPH5FmBpLvdht
gqsGfKP6Pkcj5RhOnZt1Wm1ghljNEFAc6CfE0mgVY55DfC+Q2XFwdOlNEBibBX7ODxtAJaf9QCB7
EFjkAfL+ZcDd0WVvpvaINLhlE02XCe5LMkq7tX3SdLVwfa4s44v8Q84tMuycT44+YpGbFI3wG2uo
NK3NWSX0mjlMiyQ1lU+KjSnAhHdPxLHXIlfV0tiIl1/QlMY8QqBurQ7uOv6JnhqMmI+uuc3eiIKW
6/ZAq6fyO751IeI2+Kj1xupUYb9YEyRSdBUgSt+Gy5miNQ+Gbtixx7nPBIxF9dkHWeUD1FwcCSZ3
qNrmXkj5IYkoPMGE1YcAZo0fo5ok+Pn09pvDSTwwFvNArDiFtQcAkTvT1gcsHoUeABbjLjt2Z+SC
yfIPiwILJk5IOUIWlE5RUGA/1VmqsZuRoyG4IBaRbRXL8htXcZFjcF8S8v0pAuMyoaIPxbnHNwRR
9ZvJcVc/Ju785NbfthWbEXjhb7Qeapa0FkUpDROcqQWgB/AU+xi58ugBJEC8XK3uox0Hbg4/foXV
h7oU6C/H6es/70QZmKp77BKZO85FcgqmeNzCQ7zoJpainHy+QkzplxZq5/eMIaHyqaonicXLgJ/D
/XN+uaTn8aBHmqH7mhFq28GqW4Loa5D1ROXJxPG8azKzNldyCftECYwzT4qyORcabGHn2HNU2q9C
C1qFIjgp88WI/OD87ufqGrsiaLItUOpKoxNREPMMTBI3fMnRemHwILM2hRCFXAV0uMg9X6XwmWvK
MdiCHbyzf2zHx8lw8TZgsAvZJ9mqQjcdirkiGGTDQWlf0kJOj0A2/H/OQtbZHoM7H7eLd40/+Qpv
HxekfMr1SKakTCP0Ld3waQIUdowfN7Yxg5sbjwNt6VLaovIKvf2ciuBpldY0vkSTCHS3KP0f3c1s
oo1Fr14sZ+1GaLnt+nEVtgIrXAqChEtX0MBbgq7Ex+D+4kbPY9HwbWtHJWK2yr3feH9JNqFN/f7q
aaziyaKWmXjBQU3OQEFkHQoNVKmc3t1NZtlWAoCAj8V4TiyUC8r7OvzwRZ2I+Fv9NnY3MaTPJdIC
PsX3TZhjDVn4RgCVVpUUX7PKrb9fGWhteJ70wRQVcrEktJLrxdTj6grzXjnGqXyFe0OTBQ3ERWVx
9xkq70irAMRcVuiOHxnulABBKWfaJ/qVizZwT9CgIYuqloWNC4gZ/6ZhfjGOxvUabZ3usAxO6tc2
gI1LnoACOU6piQ/F6y6X2yiF7PaexHzF1UIqp4UndjqpSZFEaUaAlgBbqWzwHwvg83vMoeLyzNof
MR3Z+gF1QC9s5j2shxC4ZhwS1cZTC8AtuCBdjdNCYuUxZ4lnGksiOkmk2BNZie20Lzn7eIGkJfVD
rE3O5hz59waI+Mo3QIT1pBb2kAES+fElsoed9YIfR/QWFZkzRkDCJMfyLhJ3iT8csYU+StBYQs5d
/hjV2ETXJNuiiJ7zpfi5mTm4RigxhyTsR4Ul6EOJuCNcqYd3HlUWrZnSPdPoapaXG2XIWHw3Hicg
OK1PIsMQ5rj0jW8p7JZoW/2ShtSSp3l167VyZjaRZo39WNq5VHOwwaSe4lDExpBHbrMxEpw+La7s
EjhRCEfiu7Xt2KeY1MElhMSEi0OBCOf6+stKzVFdCwh+FJB3UAVmMsskxleSc1l5hZgG1NnsRwCr
Ky25wMJbzvANsxmfxVbnVZDaXKzgAC6hBK8QKfa4ZT67MxbBcDZyz2mlk3clSi2WqEUZ5aoEqj67
4dd+/qS6XPWV+LNH+LIpzdyB8RL8KcF3CmWTma5ZewvVHiTdFSqT0MALd5/TO7+Wo/STpXwZPuwr
YJEGFEYw+t0rJ8Mx0oe0IwpITYeB0EaeZVn47ZLEnCxzHneIUMGDUH9/n/ZK3vqH6kgvG6KOAFMk
VD4EBmjaJR9Y3nBejUIVSdLLiW5vKC/zknx8grrFTkiayW0qx9nhkxSwMCRsCcpwfZ2hibC2917l
K2YQz+/XHv24eJ0fe61JkGOM02j5UbJCQHKT1TBVJIEzq3+0CZwcElLYP3ZhyKT7Ueugc211Sltx
Osshasfj0XLYbFHoNWzwp3wD4/T0dnJ7uzbg8wreATrE5ZnVRxZpJiWZwXPTWcjrnwLFgqfKr5Ux
cFNjxgzFi3pbYvzyN30LiXN/5mwQrZho5eeAeoIYMjRWO6XxIRhw7N8AYdheAOjx48JgolYuu0BN
GFsEqk26g38TAp8F2k9uQkPzHV6RaXswNu1EXOioJgr35aJnqgDxrUk8gz8Y2VlDl8iBlTeXLyud
NrF2Us+ggatERIBgV31a1uVytH+ZHZnMzqtjdXlxi3c8E/lAYDSHkZq+uk9m/yhOoceat/2sphCg
I3b9wlALXZjzmNmHN0Idzoz2XHLcKz4n/ojn94Y18EQIoKGsUjLr2OTfLR8CRVN3thAd08TX37Ut
BEY+jj2iX/RbCctzye+lGbqvW+ioH4TW+qgTMW+HvK5m+vHtEj+WjMqTFDuqY01uMYEbXuLR/2jT
EBzE5H6dpEC5mqdq8JJJz5Xu8lLmotRlk8w8PWpU40jOb83g//6NjI40+I2TDXBOR0gDH9CwiLvG
F1n6t6OpRk/iIE6Bw/dM3UklHakTYqv2UBbqMy3r8o2J+60EfNTXrLcVkS9Btq+xoptApc9UVtU9
GncMQiF/sxPas+AwFil0py8g4Pt2UiSHxb3T8uvgxCERgqoBk+O91RR9NAw3Trk/XMlPBksXypd6
uQb5kUz3iXxcqLa1btLAvjv8gcqBM5NDePf5Ha2B5wyzCoLWubNdQi6zaqtl3whCzexujw5OracR
TIMlAOKiIUW8nOpVB2+oy8J2fbYvPBT4mO5xF8RSCZXxIiunXgeRLNO2wF2rwmbapvQ/tcWU+Whu
/Y/2nFh9vZOMYL+7ussismuP6A+looy8etmpW5ZKTvYFpHjcHMbtxB9I6UTWCw5mqCHcDAd2Xecu
0BLuj66uLNU/jAWhY2Xm1V0bIijc6XqQCGFwpZ3m7CxlyNoxYi7wVjraFvV/QazArxAnER7aXz+s
kjUlq2zX4VlZgkTm0adg5ldfsduuRfhTcOUu+Qrsk1cyyRYT2J8h8q6lkPOfnFiqGAVKgnjUdrIA
6l9RSxiCLrZF5IaNNJhBfqcvQTh9P2YG/kp5vKXXjCDfEK5tNY59KEBIzIm5b8DV9hSaI70dVIQB
lCpFzXlrLNmp57DhCDQJHPg5occlVdknbVUpDA7iFqsKY94om4lhynAPnIpHMZ2SUMmX6eTjlqey
BybEbXbHB3yt5gw5j+vO9cu4Y+NH4beq2Er6/TgTh/GBADomyzRe67okugPG6RUlCmCSjcfSogI0
RyrorVUvOsiDVnL2Eh11EoITCDWFPhband88Kd8mkmEBe/B2ZgNOU/ZOAJhQOHibbQsmVcrkk++I
AaBw2HdOlS/x6BVLuZqmzTqz7ArqJjxeIzdW2cp3G/2pABvKv+/d3huqGcjmhkNv831C41/3jrM3
czVS8II1Pl6Gs7Ws0GWzGWpkrATB6oCt5rWyNYSl6Fpp4OmwqLvwtTQ72gjDSSHdMwIrrtUTc45D
KwO7+8icoxO2KdlhDv616qmNlhhKsQyt51IypQzoy6TX6WlVKkBOSGDJ257nnOxW/0XTWWwvip8S
457Ga9Tai00HaREZHa6n6nQxMH3W1BNZn5GQ1zJZ2EQYmyg9ehLEJvrH4HSYC9XMjmhEkNabln14
YQfyDsd6t6hwPi+LXTx6UI+URU5lhpW6Jt8gelGHJy8eeCtNtqZ9NfZY+i0GSQLx3YdvN7lclCKI
djezWStoWetIaXwwPjzZK9IzD68TxtAv4NuvhyAjhzurLuV90XZvxezcBpxF2RxF13ix/FnHkPB6
oR0ZqP8rDm2yZKkOYPG39jl8H817m0ZuNb3XVtswIPCS3Px3LBYR8WTjtILuEhC2V9JosmXvSY3Q
WcQ984DV39IFYRWCwSIPlf/BuMi45xOoF+T5q1dD2JoJ0H1AcqiBr92YUhEjiqWTkzQLxjcsmfgN
ueTHUVANs8WZ2HS9JPUYRJbBU5AKn4Sgrbg3oLeGYvJxJxCiwV8RszeFA8z0rHkxnVbW65nfMQcP
6nn+C3IYv6Hi/BHljXv10lKW4LC8ajmrbtmDYaBG4jtnsSsvGTs/iemKf7aWt4WfaOSffKP+YlO9
ZTgbljr03i5PrK+k8urr86Jwu1trHHozUrIj5vwhFOyw3BlaZmJ51B8CL6ShpA/Ayz/FVJmdIrqt
OeL4OHA6HjocvF49hy2EeHC/6YrcpqwgBm9oqzhnjLsb1U83Xxn2CXU3mqR7QSrDRyjk8SJpb1Rf
BDbCZkovCL/2o31VqBjzoHkkIPyY9V4NVocdWKHU+9mVZN1wfgOtDCjB6wjSg4tepG9JNso58hFY
aXDEn/XptzPKbHDkxM8sksKOV10X/rcwJcC/j2w2vm/5I2b5IcFP4ImYWrCBijbW+vAJ7BDjKIKs
ppeIO+87NjD3QKGYN0+DJm+3tigpoiZtoUH1cBYQiN8Z9zwAbQNIu0Xh5/wNUddSYYatm0tW9txL
Zga3QUgn3DljTR+6tUzWlvAxIK9j2/8BKSIqB0ZLuwzWVn2i90mvz2EblY+fw+zOD9TFLOVGLZVH
iv9vidfsbedjRyuxcKj9XKwy4X4s+SdqEL3+NAmQecNaFsXFnurmMEUC2fCoQkrf2mFnwTjVHIlK
IXx3fKrUV67fHsm4Ui+hBZFNNhrY/p0LxW2xSRtUPQA8YXRTBRRrFkJ/K7AYklm82MA2cBrf6qom
/v6qWQM3JpEC1Pr16X9Rb4oPtyN3XmtesFO+k1tMkKuoC+Z3L8dnO36d5AQPc9pmd2pP3rcWkuFW
QJc+D8E6qCMozt6CnPVnEo8mTGswmsvfOA9K53nwbzV9qbms5AOTXEir/GLDNyqJZ42zHVFFJgHn
4/evdtCUtsVo8uPylik/3CZuI3F1eJZOqLnhGjVVvmeOF+x+NFB3oJ8b7mVYvrZMzfZFbaE2yltj
6Hr026DwAUbd5U8pXqq3/CjMc5mYFrN4k5cadLpup0yvKwqHg2Fylkd+NGeqGjNDnB5m0FwiC8ke
hgUPsnY1w/Vjzf6e19W4cuQeBjMn9Ol6rrNAeWArtxC+0LDt9tyJrxHS12uBygluwsp9D3Lpszyc
xhJm0rRwc/QAp7L7kWr2YCGMpv+USWStCtBY7hU7wry+JYrS2hL4zXZtTHOJGmHgCiHo0Lstq9bQ
1Ym5FlFo/VurjQaOT1vjur3sXRN5uJeho2T2DJ/NPz3IBOeaFP8s9iQVUcV5MZPiy17NPktgZPb9
rnAYhui0lYdrM+umm1yTRS68yCEurWTyKH43cbzlaIipk1cow0YMqIBJbWfwE/QfApCEqZEiy94S
lz8grPtjF9kJFYw5uJr6R+AQT5j6+3Dg7W38ahu0NH6HV6LmnGKrWyjxTXgYjipTMArPckCq2c78
KPycucIKpMmtewMwGk386SRd75ZqTWAdPOy2ukklm/J38kX60XQAYExPNUaWomXWaAbx2d1rQkgr
/mUf0vH7LR8NXdm0NspNgg10nWayHMhmhuewl9FcPLzaUzkSqqAyfKIxFF1obFTWeQ5T+JliQolg
F33LbSwBeZk5crPy+WRPhKzVS26IjvZc5zjsMKYu4lvBzQfwp1PfJysJxw6U5YTe0c1FzZkayhsJ
FnDA4ZzUXJSobq9Cezpxi3MJA7JFEzPeA06SFYutM13PLMP5MbJ39RtK4u2BhxmZKrgG/5Wd5k2t
ZlKbBI1Uo7VdYCSHJ5ySzPG0tJ8D+KGnnIPLwBfOJKv+TUzuC8nnSEGeU+EYDzE+zWeJPu8eIBbQ
XobdyDbuJDau2MZmctHNDN1LRuV+1XIQoTCSk/x4mjFN3K1oYu1wzYJy6/Ayck1QTOMah4+SaXUq
LBhKG003nsuyYWtueXHIV1dSzYkeefIghpm2JdFH97n3jHC1ADR7UoaSe0dyI0biXasF510ZqumN
BeIiESoUr6m3nwpZx9GS1kIvLaqnopOUm+xqp9RK8Kok40Ao16vPgBAl1+hrMWSsLORxvlpayk8q
6S2mAAspjH1AzYbZbWs169OQm09bklaqg/ICNDx6lRDEZZVojrKNvKaWFewK2pJlQ+WpaVyk2l40
qYaqTZbfq4uerxOeY2MbKKxJSZRqTQaF6OaF0ZpuATgk7u/DN3LBg6gzDLyjplOwFnN6OAPwlfGc
YNCmagMgR1+MMF3joPAPDofavzwOGhGo4Fxniafq+KXzu4gWg8GB/mKL3draaZ4mz1juTmloArQ4
ukkRhgMqxjbNZZ/2IeOplQ2qop43+7BMrv6rdVfYHEmCBJWyW67g5x+2blOGeQTGW7O1pP40aOAs
sJDOuVd9v3T+JCTlr1VluQ+64gE15Dj8NtVQSOLrchNm1z68lbMrZsUuCTTXKwo7z/0G75osFyyL
Zi61s5sY95x0hJ6mpj+lgHuX64JX06AznFglRVVT6lnoLSaVh2teGMoyaml0EubhFAFLFSuYo5Ts
6A0tzsCTsV7br6gJ/61eK8q70awFYIF6WG4pP6P5o9U6NOPZBOnE1vRohcu8cmkk5gPSQzgShPSu
riUk8e0Fpt21G55f/rn5Ckt9lrfcCTX20hLLZodHDdIHatHHi5wrt0x76H+RNFUV80cM2Jyr6EBV
/7MT+P1nFPft2cL5ZZwj2dlo3ltIsF7aF6TrF+TZ9SuPvOf2C0Cu8VuzsufVWiVv1xSw51C4by6i
zNkrYO+2KmbOx+MgICwygfm3XL0e6+CG8ax+LJ9ig2xQwdJYqjLuiilyLWkEjTRUXChyQvuRy56L
kRefSU4XJhnrjTUICe2gVTFH+prpagtCJZi53uAFGQR5R9vQvjdYPjYM/VOr9lK/Z9RaUUluM8q5
7cv1moVkkUOCH4DDywwGFGqWBwvglIyDm36rSL1ghYKtr0LeP+5qB4ijOe6SFM/UgYBBZTFDZGeg
S3hBPekW17P3zKAP615mVfSjIP9wdayOMAnXMuH1syNirxR+QNfhVM0V5UgtE8fFwF721q7J/ucv
dd7DXM2O/9elDm5XU4dX8pxmdb1lWvowj5lgjJkDrMP0zuy/tjJEXZ8iviK0iw7eEwCYgat3SdWz
7VDvtnitAHLeJIOq0wokSE48H1zQ+DLmm1uGdl3o4ERPfC5Qv7dLuQI9F64VIPdI9cHAIOVTNao+
jOPzwdcnbWElBhJGWhZWR74psRSW+VZ+9SJ9/VS0EjNhwDEqoJWdLCKBA7zv+LQj7PI6L7bn/Yxn
Rmdj5YJ/Q4zAqBqabjDDnr2fDj8NnG8MUjuvGw2tvrZqTvr7rC0js8OLMjO7OcijZdgy3qbS/K7S
GEUuH0Vbpxy3fHosTko97ntn7FnchniHoQ04ZUcgyLtAdaGoUravnCkm0aD445lhAWqkLSC4tohT
W9Zmev5RJ31aQPA3FeaOI/PXw7xPpJm/4rsXign1bcof6vI6dpNJ13UrTpxhLhS9fcHPIHYC+Gc9
t3zLlrDsPHLTo9xhczOKo8DZD/DBQphZsU33EJwZwXcB+vaY+Q2PB3UXYLuwf2umnoWog2Vp4DQ0
fGTycTwEuw78qM/jhCi4LYxy1qfczMWwc8oGgSu6hMSdJ+X5TYz5AyNrD8molLrgclxmXsoDRAN1
vIsWoaOkMUGvHIwBLZnWzL1duGYcNEDJ5UEhq8zGgUsfwmaSmMqSFMOQsOHXL4KS8xBbUB6c1e5m
lq9WlaplbgtCIIylBJoomvP2+eLGqMepq7qfe+dyYPeBigfCMmOvOCw/H+2Yy6lDcJHU0DoVAmrP
OhlNunkOnB4XfDG95v9kY88kYIpZsFG3wY4m/ztJaop0mJ9U/gVLTW6ZEYKTUwFClf7bWb322uDN
X1lLM0lQer7cAvgUn9jLVoxCnUwFWtfxLAI3u53swR1bvOlbXMYN3XTWf45yXbPeAVfAcM1/VGFH
xkAzeRF8/KZbkTSc3al8RhXmHbG41durl5Prn5d5XBsu1NAzZLdRmu6PeFf5cdbQB5SSTgwg/Eki
BPpbBmr2afycvmeBOvznMOUUHPkOEZsgWNtlEneNnetM4NO07RppqKqxXmEKtHt8wyiA/vSzroGk
ZlUNmNb0JNdiNfVEw+k6gfXBjW/RgW6CXEHh3Z8GkM4K760MuR7d90FsBviZnyd4VBcNZCyqiOvj
cmjP3i5FsYM+ZAMaqEvu/8qK6wwj7/dkRq3kP8YfeqlOLtdEbEIVBsZv+m9s1SVfnWrxtb8W+br5
6L3Dy0UvMX9uJxCw5fug/7R/ZuhL9HshuEMaghHBSgz3Z/1bRKy7izm1GczXNyT4vOJbrrFP8zRW
jXYVlFgMh2Lde0Gki3e/JEN8lnCqFaryp6peaQCr+SKv4n2t4ZFXVEjUWI2lGX1Ib1dYvy/Z4JTs
6+AadqF6jJXzgBcKC427ikKKAnoTZ2HFB6Pwd7PUzx/waN5J+N2J8CHerE9xixrjorFDrCmAG48d
3SFVx76mw6stIvVMiaDeCmeZw7GKHFaLOSqKlstUmA1Q5RcpgjWp8oESJiOoFqxQgxKkbqnie+yv
qa/qpUf/CoICsvwQyVdBlYAsSX5YM7NlusRRw1qlozF6QOKSSE6pccFbglLNavK6lIpfafQL0YOa
aDLhsMyg5i7C2pPS8OThO3G9Do186BwK44WZvgocGsBcSI8FhaqYH3FD2EHNrYP2fIWlu6cqZOTf
GyVRDWn3qKugwMT7DenRyaMqatQCx9zy6rNNeRaDIdwGnLeHBiJ6nA5new5ieAeo3yI5r/Jr7ONU
jxGbQRf5+8L3xCFF1X8Gc42AsBYnNfupie/QvF839ZCDhc9H3HtwPTMBouGFJxoMgo1nb7N+QfKk
5wuJTmPzqiG5mTEr51FBj0BTXeLn4Ex8fCOOeA53A2WWbY8iUm/p5CvNM4G4hfkydvNxlOpI6r/B
apkTql3u/C2dsR+zS2kBynyE2+qdXS0X2V6pKStUNEt3KeNeLpU3Bm9fmxOCZAb5L9J94oWqhPVS
l7OIqZhlbArk3paSClI7oxbzFGeL0eCpp1nxhFQTSJkwiIgoOnXFAWmIPGFR+Ly+3Uv6nws7PcPU
NjJfkJKOuD2uhZURR4AG+7ivrqW/BeNMHfZrAOcOGvJOHIPFC6/XPkWq04miTgxMvpOkPT4sohNe
ipEs59FAn5ryBjchSnlcnf/azuQb7d1C7y1GGX8Tocc92117xX8MoLt2sIkmaSxp7Vc19FY4q4NO
QDjThJJDzy3nMEB9MX7k+QKQddvyg1EmRc09KnpJ9lQqShDZ38jbRWeS9WopR9EGYeLUhoQabcHW
3TpsPsmuNT+onPD8y/RSOi9DEnzz58DA666XWlBK8gYpStIZ81tFY1b4aJwrUWlLSOuMmjkShxOu
R8Lq4tP4SpvxL+UVr5h88+wMIRY46XPv/z886o4N5oADSu/HWb8VXyoLstKLTCQ9jMg+J6E/auhh
F2miIHnOQnQsyH6Te27JS4e0G9ELA2l+KkpoSjp52dmyYVl0BxQFxqrdHuHNbnJRISlmk25PjVa+
DZGMlynwrOPtTasFS2w2p/ZUWHqjN/kfIqAKg3muzkUvhdVItFJfgNOZxZfqHpLtrYB/r3mUXlXz
/151Crx5SZmFEd3weoPk2xhIJKxO0NwiaALtuqV/FJ8RiMuP1BWRCxrKo1fIEpKRSRMpybkMY+zH
wDZih19yoikPx0w72cXkRKOQ+8XfyszIR+ZL3EY/Ku0Cu4qIvXQs3rD5FA5YB+tWBNP7nYx1fMBJ
+eGxzCPlwWOqcL4Tn6YVEXe3Nk4V4wAvjey7IzCD+TcLXuhuYHoPp6D6bFeJ7wPz9lmIzNih0uSI
DbK4sRbGU/gROr1YqCx/6O6tU/Z0RDSzV6pirKb6pQa79N5YM+x7qYBNIylcnItZ8czH72ecq6GC
/moMmLz17op6xafnwfQEap8OYA5JS+5tZhLltFOkyD8zrvLqK5wzVlbD0aaIIr2f9SPMjSVxQYRS
XiVB8Js+bcfN8O3HF8acn2Rnp52icx5BJ/b8TzzU13kFSd1OESEgV++/xhzX2dxu8LrwV27qm/xU
OjarvbvBcLFXG3KgYbYAGmetD5NUCiqPaODw9Nnf41wwI2SMx1xfpugewVeRYvo+5nPzrBfOhQsu
NhqiAK9Kd/TF2/8lyEPb2cGN1GqtB5AVmPCP5Njg5x3dvqts468l650sh631Q7/FxwfrScwIQWZE
IwNKxjHBsshfJctRDH0CoHEYCbqCTD1nfjScSxya+/D19v4K1mb5CiEn/JVvAzf8aBO/hwVAMmLn
Rd0WoArGD8nRaHqnKgZuY9Rs+eYxbHk5+trFfgpdSXAga2XekS1HElPcRgEhFMZIQ5XJst4xfOsb
1Sr0nN/TrN6lmEKBJA4oirhSMlwaHSwS2wmffUJuGAj2WHveY1yGkZjWfYPWIGEP+lH3lHD8s2kB
FyAL4Q1JXtdv5aUIfkbZph2onLY9b+kPWGHR5F0UvY9Kycca1RLSIAi9TrTbBGkS9M8D04tVhoNT
0Y49m6+OkKYTQ0BW7wCzCOXD1CnhxfYhpg6PgSxAPRurpjC5Y7IPXn9XtZ+/lthAjhBoc559PCAY
qVmdfXc7B2ENK1JG78Adr2+aEhlklPrLDMVVNWfxTz3Tba7KMAZZjmPmRM1MFALBwuZr0kciX/8K
880yn5a2JY+LHM0LtcPX4EWaJ6GVh8lS1LHWwvKwR/BEHCkc/fKAMJSeHwRmp7V/K/sjujPIPqOG
0R/G8M9PH30uS3ZWX4sDSeMbg7LanJbVjaAxtyoSSETxehCE8OJX6qTJ00DF2vlDivlyBpjti428
5Ae0FHADQ35Q+h5HV9temdP4pVKXIbWwBgjfUF1FtSyvtu8N4HSaP0CCJwVTdWD8xkCwUJDIkZAI
C1M65Nl4wGEHX2aw8x+nVnFHZdJGRtm/owVd/V42gZ5AnpSB/OsUxMHBK0MjBDsJ/uTZ4l1p3RKR
0fJcvDDT98s5N3TVQTO0BydAtgMBNKJb8UADdXteTPsrh6G1yE7v791UkLADnHzNTejQChEuffwv
G5Rn1/ZwQZw+ScU0Qoajaa7GLX+0vP018caF0CGhxqCLO+IW/elqJMfxnuHo4wxmCyUU6uFjbnzh
vRwPy8QS1IZF7dN50ipiXwrvqrWeiFdtqko+FZqj5M36Lb+rqx8AXf3FnuIePdy2AZb9x0AtJ4St
I4EthsH/AT3y4pYinkTCBXgkwgOO7ICp23Fk5eMvmTXIsSVz9KL85obky2ulXxCX5vYLOWjD4TQs
NpJ/QBznWXuAH7fdmZ4WDou9PpONbOgfoIk/n5xuRsO1sxmDdKHio/nsIfqkM9tNpCbFrdPg3FVl
WRQwkDg2JuivBeqCVo1XLNJYlv4kulzNAq+pb4b9nfCtk+r2HkbB4+HX+gD/h1kPhn3D/jey9cPg
W7wRoGrnIChBAM6RG3ZdAb5qLx5nzphAaiHpUGq5G71lyW8xrjE+fhm5OjacSEGo+5UfR73uDUmM
4YFuSltZMiIbkaVzgXzHI+piXb9CqN4tujLPS6R74S5biVsl4wNG/umf4X1GkiT30lm40AUWCJfD
2XXmIvc3KbpEnx4bphmK0/0Lx7F8DmiNGAZ6o8R7ob2os1+7NCKDePgqnawI84i2uqWTNf60e+l+
wrJt0VZJudO/AU/LX1tNyIwDGwrDXMyXDRxcM7ogsPZCmdtCUc/v2R9YrdAXjT2OwSP1TfklMcfA
cFlc/p1XidUW/Taeo2yOWtYOZZug9NvbFMhLC7cKJbLuQLz7GX/2I19Sn9IoTC+zI7jBydvjmPvm
a6ZOaadpNE5+PvSMLu7HQthp14sIJFy8DHKb2rTMt88ttOLuhBjbf6GvPdN47a5+GjDw7d1Jh8H7
6d8FdpzD7eHD35G3x+Ms/QToGwovgCtUscT4ii3PUX8nLZjopxB0k16TomvDtWmDYJkSJapQEBPd
Z/FMOFpBxqqmVbj17HBD8zLmptgI9fyR9KLFMw+PBOO+SP4q9zrA5EKK+tqowJQbbEMBJ5r+fBAm
4yo8m5RV8bJrwRmSIUUwXgNn18DpnW7C5g6Ch4lsEseBh5NLdZQgHCXPXtCp8F1uHZOmBWkpLIe7
YagmvyuKA/Qem3mqUCdRn0yAMHFBmOGePvK2VT5bo7xkKAdObWty8+SMjrYHkagGanlxXd4t0XRZ
/aryNdAfdncIaFMWfcgb+qzPeOBvbItO+WsZaWIpXOe3nwkUK7y4ftJj/wcRoYzh3+0Wvpf2co/y
UdEqKiDGa3E6ya1ZKra5dZpk9b4RWcpuauBRHBUt2qO32ixPKHTxTvaZj8bidR3Yzjt+4AXCEXkR
DcHMVl8rnTDUFLjtzdz1uaGoyizT6eKEPrAdA/DcWFuZeWdLi1SOCdPgsMEeuDM40SYAKotXAbES
uw+xxRoGobwjWt+3+5O04UBuB/ExhIOec/8/BULXALvnKnVFR8TfeQaJ0XzXHdxFeX1RjzvnGDXT
dTkxV83VQ4aDLVgJwTen6bdQvREGnNy1rD+YLmlPlY1AyORlG7GEj66g+oRo8IoVm6hwZbfylLUx
yPJcAgdObmbHH/KiXz9591o6YicH4OH64UGuNS+UwtVmNV55eXz6X9/Fp7PdYmf3xrz4uJJEAU67
e+doXXkOGYJsKnM0PJkalH8zjf41ohqzOS8MxTrzrnTiiD7oQyQspW0o7KsAZH8lP0VL03WuaVBT
BxFZ8kOWyuEC+EE2GN1BDrfnTpTiwGttat2Ew1tv/lcqhmY7z6uNREB5LRSOOI17Bm1hsFwO8mdu
vcB1CvXAbkvjwvoUsHop1cXAvVqUa4b5I7eDGMqeIvx1lVD21HIBNeY17ulYJpQpB9SVbmrpC5jC
rFlyeBdh7dG08oMJq9bIuFOttYkJrvNCDnzE30svg7TTkDABKunQ3s1Na/gNy9Mkq0yFGvxtJdIY
juGo5P2nSf2q1aets1RPstcSr1gjScSxKvkzYcZizzIvRDkq/fSkD8QoxlOOMjQyeAMcTBVOqCHt
zJ8WwBl/os2/8ZEaSE6y5RNPc31+dUSto8SMEXNNYJYbembvUSysMs3hQyuuj70+W5y3Lz5FYNjR
I58on3Fhrjs+wRBw8KLvFeBMT+1dfDjd0xGoVDvCe6v2oUiG0kXdFxalX4v/ZDfyymCwl739031Q
RsyR8qjbWzD/17rHt7o1955m2PnTviaqVLeeBY1zC0TPu4Q+6SDG3kc0SV3F4h1SCse2VqIPXivg
uqLq+UBPFlbag645FNQnh4mmuf4OcFM6I6H/G5VtSbsV++XIrXeuL1xFWpNkhF2GjHKbxKFWpdka
LJs0ZWoMnDRFDqYjit2h7uRtlyCurPww0Epnl/6aBFLaGieV5qo6DtwIRcml4ElSyolQsqcXcW73
bYchjnlyadrE65Vc4qd7K2D35NwjVNAYSbYY/c4aEgd6nnVSXeExotfria7pAVIUhQK5KrFwI0sP
jRmMoBeKUThwp/huGnvNdVHFb48Qs5yEC8aJ1l3rIQx6oiifkIxYR1xoyBdtQEhIuuVBYK/DHHEt
NHa0VNfoRClLNEybEuuepqoTHuabA1xBXwb3OUZW3Fhv+6WlBf7noCh6rhNmejK3mvFNb1AjxTXp
keruGCC5x1LUHsl9tOywT47G6amiV/CC6R/4E6G4zMa6Ju5hBN806go4imu1ktS7CZOPatNowueD
H4Ss8WzpmPas4yWk9uD0wzSYwlIjjkE3Xza244dM/BnUUmhEoAa2V5i+ew1lv//NKTyxl1ixIwsm
TNUNuM3k7T9Jl1LH3Q/N3TSnpzYzcMvTL4UuCRUB5Iw+UtETWvExI+kca0lC7lCnMFBpoYuPNOuO
Kl25xoD2z+lXXJ7JFqUqka7sXUcvWNYzjVxDoMvEulnAnqEApiPRPx8Re4XsyXLktJ+wfc6lO4Q5
wDpqZ/bIEyu17W45BVbcEeWweMLKZBvKb8ic74lz7HdukWnqAJQle78hGPO9nvrHcbNnZcz/kuQs
5rf+g2hs+g0a5U50q39Tbu/HiqXdet5GH6OdQS+XcnDEaGoLr61AohwHMOMg27Co6OxCBeJmQpJb
WwoXiXV92Hu4679lHtTr4YaZxAf8cdPZZucryY4h57nQyRv/+VGFVJgTWBttbsdvv9jRmRHXXJ8j
K13Oo8qRt5+64HtRVZJv5d9z84m68ptfWOoYvoNImB7lr3ncw91wqgwB2IortQdFiiLJvlA41t28
+kxIXZGVvUpMIuE+4JDH0LjeLA2oAFMDJ/xqJWUOT/X8Jn6rJh8e2ZznXqQVkpNMjVQ+GMvVyETA
JHo+SivVwrE0n/YuYiYOSk8TXCu8+aOvlfuktpV1CDomxCy3S0WBbLvps2TCsVdOfyMwDOOlqJUF
Y5mKtkFGjXtd7ATtM1pAj/7taDd0EpwxvXkUaf5dm0El68QBhAngjIdqAMWZpDOQ0rDU51qah3ep
KN5O64hELCBg+h1atymE9Nvw53Pbja5Bz0WPbpE4XvWMKpN70Qm97G65oWOVzbuKOnsZAX+0e1zE
bnCpk3AcKpp/Y7uA5dVyY7lR66P/5aAqElsV9NliNLogETq6nVdfHmt45JIpEQoNnj+4TG/pK2P8
Gef+3O6Ttm0wmDL1iLQTE+PY0f7gYHKvvqIwqkUXiPmul7CnXy4XZ/uSEb98qt32tyNZP2ZQOs3M
+JHnKZK+9ir/SxmltkexQGVw2ESyQOEk+7y2kMngKVR6fspsKkDAW3eKVVYN1WOB6Rm8f8lI7NHw
NVdNTRbv4zuFBhdrunzeX5mEJ/yjzgF5brSttht1ZDEuivcGZTNcQDIH1GMWCB6Fml2cV0nDur7D
ZseZHwiDLFDcEaac/TVcYMogx3GqNAn1Z68VNug+3Nwz0aGPpdLusvbnBcfRyapQSMBDVHsw5rwd
oBdk9ROEUp2K4oWZS6C3pii1Mcz/689h74/6ump5xFkThwfOPp/BjrJD7yAOptDJQGCQeKQH7X0B
mP8Ih2RBGYUJIRK2ZSYBrOnZuR2yhk8TepxgQGv8HaFsguv/y4v1BgpI5UuLw7RanHKN5kndC8V1
coQrIA1oaYFo5GgYalwHNj9AzviMFAU1EnFukQWZzwDdXUrT3OHTTXZFuqFbnpIDWq4gYgA+N96Z
GSiuVLZsNjqZeUTH9JrtoA1ZeymJwSPgzfZBUoY+mKeDnXmpoWuXpmVK0y4g6dyt+aI0HrBfejQx
5L/zAoQRdki2gP0UjFh7JFRe9Q2jnKhgI1c+PhOCy9mQJdX2nJsN43i3d0Ljh38kBdoklX0nhVg1
1ArExQOjKPTKlAww3/iwZueYRddCOQdfgAusmr2lRGNqg/Y9kBZZED5DC9Ho6flZNo7YrkDWXt6H
UL6l+olc1IjyBsMZS+3Sp7lN6TiM4sGQJx63axXU6tI+KwfCPl1FFzerVJwdNMqPpQMfMkiX7Der
NGZWTnvWBw/oHPE8ug/KZAVJ8eaFr9gaR8FXLvg9TNSxhwnwg9Ev5C2QmKiVVSQjwdrvfPu8Ft3y
3bvTt3k9oclTiFgdTYwM8Qh1IkTD+11RxrSYWLWQlX5M+WM2zkRTlvakRmXtb2hJ9XE4OkUqCu6M
2OSW1fTUItp197Sk2YzSnLNNsojo873uk2pd4kLY8rhLXGpTTM0iqbgLSUaF498gyYXA4TmJrycz
FYL9GLLqSTJjwBpl1QPfCvk0k2JRtWjk6KmebTqkwpkZcMGQnazXCQgbGih5kXaGlPXkOExaslCs
PszjbZiZ9dYQVyaJfWBjZ5M/9bPCX50hw4Hga3hSj9Ynwt24EFLmUZwIm411TyLnmFIBwz+dL7Ac
Z021ZypbcBfGBJESqWRMUwQSu4eDXyVdELiU/ZfIHHmH/S6jrXtlfDBumMINnrOGrqlDAl+qsY3E
2RyeEWZJzSRjSM6njaraJV5ByUXWZjppul9H8nkcQN2TjfWEFq07kcMSbA0e2PurAqg687dybwop
3e6eyQ/y/0drq/8gBvYvHJSzFWjvC1kY+3+aQYu+XTsGH1I20taX96gVS0UmQKAFCP7gunieuuVl
hkoO6rO7y8BUqAxKweByWAx6kWrjzjO6/m03+OGRkshgL248HfrHNmt4Q5yHZB1T9cAEsqcIPPYb
cc0JtwTPo60zybMhK6bcXSkOOz0ahI168YD8VgUVTwxjtvcBcTVyJNB6qDVDXSVOzdC2gOSifFgB
UCJviwIz9oWuVUkJPWtKWW/S7YnbHFFcZ/rgqPobBZWLXIVUab242rzBqHM1HrfozF0iTjt9MfMn
KWCrRr7qwgP5XoeLTM3bvoM4x4rdLbDRh+IhZu5Mz8Qlf6WTh0M46Bsf5/dyihSr3vRwlnmYsj2O
PUkW+Bw6Ag6Lg+uYYNdSFLi2QDDJQ6mKeX868Talz4YYKiHoONMkzkaInucT69mAuJLiA7ITRsNy
KBIr+Nyf97XT2nOSBXRAnYUgiFj3KPNckUXa5y8cPsIxB16J67tYMgabKVYCQw+TaYzT23eeam4u
mzX3OUbY5IU5yvaL/wGLfM/pxhpFE8iyj19j6AuGvyjCatgzv+adbm8CmfQ3h64D9dgTW+zj+N68
CUSSlik7kwnSda++ywfH5kqQ9IdbnU4FqZ8tkeudkTJu7Jl76ikvU1kVVVJ0o/QD8vc9Jji9H8/o
2Cp64BpmmvVzu98Ps+5FHa4DjX3Bbvy8/d6ZuTrgVC9OtL20GqVwOLZB1Dr3a3F6eOQ/M2tsXOnG
jZpxUwI91srR+CXQ7eCQHWV+pyaGSp6G6SjXovqWXPEfNc9qopA46cEZRH13sAaWhYfVNe70ZF2a
veKJCnkghXce3bstd8jPbOJ24nRRQk7Hbf+4ITXPnaEaXEMBR0YdBm0TgV0nwW799f1xfMwXkCKU
aeelKmjCDNJeS9xe04S+wP/7/SLz86JYJGBVmZSx5VoK/1pXkUoxvYTj15w9vSbufket/dkHFCbe
gd+Wv4RbMGA1mfe9UilpmWeEyAzHxRpz67H2SYPlT4W9fqFlbamK07C5uYGFxSu81ezDXmv9TEg9
gHrgrDrl8RjWN5aeZlGr+tpOGBL+V9M+gLqTT09YDMSiPyrBpDmxEJ2snggCRnHrmW38sINsp9Jf
i32u9qsbubZtyA4GKOY33ulJldCIWVbHhWveEMF/ICIuirXRypLfd7lxJuTA+5wg77m13GlouL+p
rnJuY0Q/OxDX7p+y7eTmHOY0q2AnRoTo8IRXixNHxWr7xKSI4k9DKcupwJZsr8SkiVUzYQZ9v9cp
zcH9QYLiodpj306kSjmRCv1TYx0RLvO0EIfzROEoZa95qrpcD13ZkPg36e/VC8RlNKUa3+ToI6d2
79zOm+ikR7zZsXY1JFXiujkeQEBMWy0XH/71TxiKKiUcMEhe4lcNdecnnOFXZZWshcAMlOQGZWc9
pfeXXbmP8PyqZ85hQtOsIfNj7HsQN12IrqzB24jKwP/m+RFx5nxX7IfYksDLNMUc1t/Sq5oOT0B5
hhgkHrK/lDHZpsXYeLqGNHWuP+WucS2rwopve9FwNH8nnj5h2Hy9THzwz7m1oO8oUxe9h6z2Iyby
29dnStub/pfSOFfWpxpN1USH+rPh2cxtyYMUiFeu80ClIFLOvj/fK5B9bw2QL83x3h0QpFeKOIL0
pq3dNZPJ3FFMvpLmplRhF1cHJRS97mr5KUGk2q5WCLQnIUjstYpt5b2nNledi6axPr2TDJv9Mh+D
OG/lh7hn+YakFW/MLfjcp3y6jK3K5u+Qp7g7cYOP1BZIQ20SFYlj5HRv/i4DNX5+0l5rztIzWTw5
5Hx0JH18cCiPxWlU4VtNTrGF520sNgxs3VvayndkZDgSbPOcK/2Kh2qrGA6rp5FGomGNMZYxj5LS
qz2L432DRrQH5+IF474uRI2X6NWjiQ2Vh/oCT+Uz+HAk7MQ1v9RWp9UWRtwOC0COiLYF+FQJqVcB
428K9jAyZz2yFt3+8lobLyCFLvDxLr9acY79szHIOE0REZ90ciAkBFlelgwuzQ0TS0CwYzDyaVIo
hwCQsuB3Hnozmuc92o//UAT5QqQRyZS8oXBhkAzQTZLhJcFWT2VrU6LfTbP6dB0f6UJ5oWSXL3SM
z68Qh38fm/Lcz2BBkSUzsZr2TqGrWVwgD7UGFsgRrRQUBIoTdhvVQvpD9PucRW3OjCOTwSWLYTHL
UTzx24A8lJe2/wo7jV2g0gaAQP5M1HIZd2LotPPopl6wQSHDXuelsNNct7X+jXy/lHR7pcxbn1ob
Bt6ZMC3MiYR2l8+hoiQJUYSn7siuI/5SkejUzpMHO1d/16X31MmzfEdy+dDkIH6YFCEEGExNrOmK
gM17tjVaY2FHl/QP0FYGxeF9w6nu73unIBa4il8LHICp1hb8SHrJCai/HwqlhbhEB4jdA6lIiCnA
btvdwOByz/VmRFUrPdrYuKXmLbj2Q7OCEAlPqoFDTK4yPcWwqD33N8WQPV3CNebLU/LxXKogOn+2
hTjQk1F3/GzEaQ9cD1w/PpRaIH3iW/j8QY5c5lB48cVmYO5Dpr4cqSD+T0E+zR2sXaW3Y770LU9t
XFilv0/+ix3b46ZSgF0EX4FGZxv+VxsjVpRuap89iNmwoHT3GKgJp05dJkJEdvOvqOL3vP9fqfhc
G1uSdvlA8tneMx/ArHXkb31sLMjQE6EfuSvZISYfqFp4qkp3HgS4KrFCyrdZmjY7bw9ic9B1tEVm
PGBft4Ul7XuJlaBRJl1/gqmLKxzPUBdN52CEFefWriKqfpvq3SyQH5i4A9yyv9j7hDrSLIpz3d4O
K0tAik452DiB8TkwNs1RudeoopMxuMwEsGUd4CALjQiLdFqfjNPFgc0znH7l14YpLEd3CckWBizL
VIEebCBJD2SF1r7WRwlOSfGR4h8BWPvtHQ6HWWiQbUChA3WukUnN9XwD7H3sfkP4pWR14cdFcG7C
a22rbWREEH3QfPEGHtBkoZ4AcAKd/F6J+yP4e4efe9EEtiR8dYezQVrBI02SNAFP3B/7V72xtAxm
74ab6z7HLOWHoZRAq7d2Wv/vFKHu3PzVEoE1C8vQYvcmSGqB5vewXMWBS3Q2b8JimhcRGMjLpjdu
14M2R3EgVGJ445F018HGXoZKKCIWlhJCCTkurLbygmE6AkpP0N1yUu7cttQz7AF3MEMEFYIPk/AA
m9KaXkcyYo/RSFqXkqAH5ax1Zy+OfemIXqjVGeI+EgVJMqKVe8S6XGSofgR+hnrmwO0WIVui0037
YwYgqYi+5+qwhGO7SMkicbKnSGhKHzkqP4qRJUeliFOkmIWLGQfklDpJmwS5pgFXGg49zRcBbyLb
nvGu83y7U0VBWcLYK2WrOPgG0D4hlWzW/aBSdt6cSf6xFX0w5CrWkdHu4pwG+a/JFoZcWsHr5CV+
O5+yEMzBtuNhGqcod+PvS9fo5sNf185IP1QOrYvjKqbq3IZdzsHW5mfORdplmyHQfziuNjPWz+DG
5h5BZTztu+c0/8Q7apAsMb/2c/1rho72z7I0Eiechim3lm/CpINLIyZvmKZgU1uyCDB/uBF0rjmX
DDQsdLU61PEkSDEvMqRC2xlUZ9nbEdWVpEY1y2ClvT8LFRK62KuyLotMEo1ummTm8xoVdkkBxy0V
QP5jF96flGmmPg7wSkXE9ppr4lygPA5T1c9ONJwt83kQRdiFbJsnhLTqp6tuTkk5x6I91/a1UPpd
/e5IVpuZEshobrTvMEJJmdiH5aQHHqw3Q0aEzw24CkvVv/i0CjRdL4tzjBQkIbseqjUaNN35H3k6
0vOP+gwLRqylGoTmCcY0JFxlSQ7fNEyGhzrCIaZP8b5QlbIFH1oBgAKS5If5zgutHFp6az/y0pDd
9M55C/SGmxBRlBumQFjh6Hmkg702corSkbQuGmKYC3PAHZ4sModJFsDgj670GqxeQBPk8dogwI2F
DcRd8uZqidDl5z9auvNKcKgYIn5CT9NyZ6V4pQSSj+6jhtZYGzPaZqcjpFYWeGcHmb5VVZ6okArQ
qcRIL34cY0/LAw7RSl+WsN2bOh+vtg6DPJynV3ulwOVWU/gXf7PdR6nyuMFjFWDJvc6gmha/d0M6
yLQCFXUcrNFncJVL5rAvAIQ9ghVtWu31VbeqJZp+Atapb+CLW8zRU2571rwfr2Jrf6sszj9Gbp+v
jKvvTTtTAMXby9BSCwRS9dAU1HXV/ma0UORlmKpc2edEBS3RZaHRQdT4t+K9wov+ouNJckdOY67g
U/FcW917M9qhX2SCiOOssvxG4XgNdExUrrptMjOAq/1RO9uwTCZip5/0omjsySYMJoXR/iW2SUI8
1+PPb3FP5pCY+WCsJqWRPNK8AYZ/4hqSst8m8b5pAWul+pPFwNC1X3erKzHu1SVcXGgL6XJcAC2e
U3CBbLE1LH7GbEyji746W3gw+3EUSUsoSFR284RRqlhhDO0LIv+rF2EyCijPkwYxwI+4CILoumqo
9i6vcrVWja+/qU64MBG7SNjwL1B0unuelyOgOgCjvH5MY6mqWGU64JqTGJNwrE4TOuFrvSCgo+gB
/8ajrGYOeEfPrucCyTx6E6YL/nL7qrLcSLk2WDX1pBezSQYjpPL7hWSaYMobSJ9ERh+XWxQyFIFt
CCH/I6j9XsuuMQdZEpTpd8NISctg+bNpZ9JUv0WFc4Jy7UOB5rPbx55txuTUK60IV5WVe8B+ZYHN
pSFu2S3/oJxeNFSas9qOQbJ83MRoWnyxXUSy7wm874/HAUaBAZCO9Fikbpi8EH62CJaLLPitnxKT
9GNcTshAvPdialNkXC4VOvKuFQgdDVIOA4RcwPpoYdb9Qd0FJrw0cx+7quUl5rm/L3KN4MBOPnC/
1W5V2Mrwol4Ifj9m6yRHx4xagg5ilfSTjZ8YwC+95TVEUntpFbrMGdiOnhoJJcDEGjp/o4R/3Gp3
8NvMC3LTp1cOzGXMf5JHg/2vBsuV13n7gyGC8hs8aCaC2xof/R+okIUlkskVxPoFAOe1gwX0MHqc
4eNNglB60/70McC854pAv8ZB3Q04y+SHPYsHiXC1UNK8wFOzN57/h7efRGhLyd/ANzXyho6ra9dE
ftgj1hmpaqNVnk7DIThnASMYJrlCgSmpJ7dRxD/Q2mKkXPKWDkcv0TZvYMrO69WEqYKHGAkVEOKC
6IfcYWBv/e0bBDkuiBBQSlBnjKIPkBxZ/P57QNyM09HKldddZbsbBioGpHxegDRIcVxm0+SHwyOj
MJBmew+AA9/qKwnLUKKxUSOh/uVnGSsXhjtTmiWt/A4wHRICqaRz7zhRHtSFR5HMq/ymVG5oai3G
M75BZ00MP+ayi/APqoTgnQM5ugHiuSNqZ+aOhp9yl96dFitc0FR+Fw6JjKwUMtfRLLFZnbSB0a5B
gUAen/jmvFaYnVJJTPPadD3ZB395eGa6RNMqoMXXXwraHPNVkAF6ojYzDqqT/OVWb6QR2unIKrNh
xeQshARulu0WBt9PW8oTdWtQwIA/K5bJ6PiO+jm4A+FsBTQeAFNuCIbXrTfujECCZ7ho1sCsi+iS
3qy84s71aUJmhppNiYkV+u/9J+T5pUjMoHYhdn77BZ6s3KtBzx6Xr8Q4dquSJUP2dun+1ke3xWd7
Sf0j58OZKc2qfpdeK2vW8z8Eac1DELi2wI6hT3heYyn7thF6Iuc0hiyAXRWYq9VCmFLiJAS749zW
aAAlvn9fCRERoQzbEbBEfMKzGHxg3FRBNwdPpqXL+qswS+TVtETNO1JZmoaTgkMm39Qga0VkJE7k
Vc8/XkzmCXjeWWW580QJw8cWaddr+LX0QQO1xAanWRJVSDmcYZXKeHcJbMkXD/v/JS6cTDh30x5B
GewY3mbwk26xQU78rLABx+u0DLCrLyGpK2+F1UDgLU+/4kIZ0l8anjOx9WZf+m8qC4pUvU+nzAtA
v/rm6y4XbXHa+KS0s7JnpF1ekyuldzstOtud15AfWTiLHma/AflHhQ0Y47NNEZ1JGu0fQb+Iye3k
nbdMaTTmp7Lapyyxr0SaSgm11glxKn8z5NXi7v+eCIXFt1qaQmf6Mhw5U4irNkkaJpVaYgL21Cuy
/aP4+1sog/GEGBE2YQrS/3+UgMEsfmJp/LSGIjlQ2wddnFawG4s2Wn2uVNdcBUmHMxzAoOi55GM4
vQ1N76Tju6m6I6c7DZv8ep16PTF3yCfesvOfrWT9HVXAAiCDC0ey34kv057IMQCIqDv52TrDxP/2
P8SunUAeqRlfccdvQLqPIOcr0nCknLuJaE9VpdCX6yOnHpryko46p0WGIyfGJa08FcinYPEvjXFb
NmX3DIrjXuYsJHj5YbhXJG+aK5ynB6HAX8NGCClW67/A4zcMYN9m3SJgmZzd0gy88D5kRLvDUfAT
i6tlHgkGe9mpbLS46AHQw8SOTH9hxurkDKAROwy4jGgKhd0ThIckQ1W2eM17/IvIMYizuXDCIp/l
jbG5kFwa+1BjuILl1azFqgYcNqr9TSZ8rSSGK07q4uYr0/GoSKydTs09F4mfE/D9pVMCcGqZxVVd
bHeo+xE7hNNeZ3QemILfYlmSCuhZJrh8qm2TL0DwhWO7ly0FRJioL+73/UX4QEKjI3BhQX7OFJV4
7HXpM6qsh1UDCqK/H2zg7+MLH+zWjahwPCcEND577Eze5nKhgvPXJts8BH6/4jtBiYK9hX/ww4KO
mLXU7Cg/9/BBHrk+wQ71+gq6iSI+rQO/nMMDXec2dz4vqcidKei1EUiJyPxT1ANzPgl69nz98kD5
WL4E/NcPz9zsJga4ih+cOW02XsFiT+EkASOL9vjcaVUkYKbcwYczjnRzVhID1umIgry49MySS7ws
RHqpeqWhXqFRZwvS9F+eK9BU2HOzRuEaQS+dOr46idgVSYNKktMMguh8Ldq5KYYq0qqbdsqrPq3c
X7huDT+Rp42gZZRGg4iZ5KFf45RjEdhSQYJnQEXSOOHGAorXrJDmjNP7yu3DHhNwoioOdq5NUuYP
gxtfs1z7+TGrRMypbqGGohfXJy2B5I/f8Hs30fGrp8k0X847CphwaWji+YrONSNJxYBsyUv+dfRA
wGnr9q1BUm4dSHdu6e19tOzoIVULofETPupejXbzOLChBCBH5dzR367IbTiRziP+XfME4bKRYQxW
HtIwljVq6AA9LoYSgA6r2KcvjLRZVwik2y0MZACqXI/8DA47TRN9EUwBaTbw1V9cM3LbmiE70Fgo
po22/ASJ0/aQfxxJvEUQqX9Ue9ao9UdyZZNBeM7M9iFGjeolodm+Dm3r4+Yh99QUUu7R4dZkqULH
gZaxmsL8W95NVoqGMSW3HC2gxM3Uoar2C3GXrAFyZcDdewZe056DiI+uulNMUYtQ7lpGX5+7qEZ8
pw83P6pKQBFF+v7l8HihoOnYHakeRsWhTD0YP+UEIovuDUmf87utf/i8ZDE0Hmw040K+FpviolKn
YjMaw4OGbiAbG7EkyPqvZ7P8hGCcjRqJmQJDtHyKBYqzey5g3XCBVh0+epPxC+Fu5faW650Wr7BG
lPBKuIhpFAuGFqvHrRJ6lL29a9WISVpieNL+aZmaCcrmqZlNlaG51Fe61HmWpimbzpmolx/tj2ca
Db0N/eqVtBPmGT307T5hfaG7fSkCWra/WPhTmM9Khn30ZGOmdixU25H8q/l9R9PPYTWU0ezEL4Pz
NyIc1GfN6ZQbahLjRpXbTzcM5iciIdxm7WKrn7YIfYldrjkQB6wEiQALBYAXssZPGvDuPlB0m1jV
79z8yq4HPeHO+XO0w5EIXO84Ia0lNyUhTcdV8sAlFIRtdfNEYZEVUB6OZKash/y787OCsXcIwH83
6KxtdMcWx1UhM5ETIA6F9BOvPvtUHitwjD/uf2peO/GXMuUj3mttmCGMDG4CHcXsDE7KZCZWB68K
jUgEXLbTd/XYnE2oDyu3N2/QLe9HetVHQVR8jfwVVpWmgOMupgL5H6cA0XbTWVu1ku9sYd1yTeEE
9CoWGtnYwv6u6KImPGUSTbJKiod6SyNsydnRQ7f3z5NXQ0pt0p+dpP6vn0XfPU10MKSc+yyWj0b0
kqX1uJxSZKgVsiLeQyHN8WEyWgNt3wsO6CYluicVy7PSqerTZvQheDu6t1pMu2Dz51/aAofRsjCz
HFG2Hw58uyXf4Au6TmZOzOoFAk7Xl+bQYM4+y8apPUyZh/YK+sU+WFZa1D8qOqAEncQZ/MdmQjk+
HhjET1HdsWqHj7Ae3wwXNvBv4YwnQhTtMNjBkebTdWvyqfXQnE5Xmx6sSX/8pJ+h9Dw/mPMfKjBg
ie/iq38yc13mNoOH8L9A1a1h/UpcopONR1tLlwyL6hMjTlxb3k69b+Xsvk15Lhge5EAzSHX9+skg
yt+Cg9O6Jz0/ShtNZP+ZLD0R2pqv5GClUJ7GsZvy2+JKUkGg+kpAEijSuLLunNBtYgIGe4G6hjRy
nsCpxT5sW+JAUT+GSjtdMHpCDrWE+r3LYLERp5va3ao9lbJx8mLn0Xm+4wFJaNWWdTtKN6TtH5g5
m3/imgbyLbjtF5uBea2ccwRzjQ71+zzKC3z9sKpn5kKGOcaVFCgTFnNu2urpXRNZgm0foxYRDcaa
5Uo4h9TlifhXuwghp1wFe9SJN9VZVy1DhwWMVDxSkKX25WkzxKJf+kif2VH1wYxXGFh5N60yv+fz
7Ff7HB2w74JzDkGRtaAfs//O5nX+tV5ZO9l5dwPlr9EF8uE5Y6iZQbtHcKsbU+7Wb/Vp2pXI8QdF
fD5un5F4E8uhdKeg3Pl2RGhVzEQ9KHDlAWwv5cTtrjRPpX95dkDV9wO0fudHMqNsTkkgqMnxT6DV
Qhrs8ITLlx/JPxg9JOOZJLXu52oyXo0Ovo2kfMFqHJicrPkYJ/WZzhMHx4T8IBMA30y5/w9AH90y
tvPLYod6YrxAsi5MaCSjdqxNfZrKgK1KytN486wQ0LRPMKhvS2xrtU9A2JAEL4t52N79dEKJRXEc
RFEx5MG2j0qcFSjvbEiGm5i3UYTQKzZjRKBC8OG+NM5U+jbYewshC+kKrWJYGXXGABE0dQ1Luwhr
CBInAiXfzOFL0IIsPuH6iafuKfnOWnFr2KTIdBCBF08F56ONxWif+CNMROLbHWZP8FZp83SWEdjr
YSXAofbUOuY28nAMZ8tyIBoza1OVjyGSyQHF/Pnxort3CrCKwrzJgnsqW+qxR3X5Y/wV06YIMitD
etMVRDuKMa0fBw+aakL3FaFhqyEgp+A0NZFwJEUGIxxt/7qdDjL2GVkwL9Kpt3JHmniQtzBk6Ol8
pGjpBQ3KAv7UFLrCSwqVkXsR+NoMJfAJToBJugvZkBQ48ukEYbaSIRuSH7qGXb7RzOpiwkslswGB
wz/GMWYvIxutQuXimSF6brDQRccA9iuldnAiSYBy0/8a03Z+YF/K8VeSmJ7qZI/psgtIkxV92uS1
wIwW/Qd59Vr1686d6QNoBBmuKr+9tW1G29bkNMxl0vcNIAuUV0jUfe6+Wgg1Rmlkf+Dr0H57mUDP
5bOUyLhyu6y1NGyKNiNa5MOLzcLX14B7x2y41cobggfWYrtxyL5oxCh38SrkoP35IybRlmGmNWGb
uYXpYWXtH1AUuxeJvI5VFoooKcnCfIHZLyXN6OG3nuPzyM6QC+9tkUYEeBEgiJWA7AnuFm4ID4H+
IrjV1zhKK2wCVvPOL1hdlWIMoD5KJDYLEQ+BTWgMMRRE93G86JSkVBPlh8sMcx9Ak2A95Rawl9g1
N08e3x/lv5MCg2Jj2m5cob3uomMNOGucVMs/ekIRy3w3OXqyDfFG81pGwjkVH+gYCIVxBJnaCnmW
XkZ5iPmm95roA7mrwcJ26QR+9G+WVnLJyYpEyEHbErh/FM39qT1qCWvULWWpZypO0BF5XTaIe+v/
/l5ZjDBON3WcPq/YhM+dVx9YZAwK6PmgLotjy7A8nPfF6cpYdJdMDR1xUM7qXQa2S+h3Wgh4fUsL
iJeJFKPQmzEs8f+79JJt+FdVn4be76yirzSpA4L9V31aM65MKWP64+2yuBw8iijWW0+owEv+EjOa
t9S5ZrTUgrvEMYIcKJ8k24oB9VvtNrdizwDMLhbNzV83d7WkZN5p+jClDPjZVf5ZDOk3eaKEwyrd
A9OrJ0yYp8buMRoJXfDG39rlX0iQfGhI6HdoRPtvprxJ5rtxZBJ6U5jjFMSXVM4CYRCaBmHKWiIH
PDieNBN13+xR4VKB2py4dSRb7N+2Vg3DiHJ1bjcMzIl5NdAOBpRjpP3FNHl9eXRbG9LP4H4xukc/
Snm7bjB9c47VN6yDbM4V85dY+2G/ZsNHh2tTMW2l8ZSmxJWItPs8g/Zujc/noaxNX3bgwny5wMEB
+i+4OSX7qzgDVJTxCB3G90ItWj+D/84UNHf8oVC7CO5M5e71do+Xps2aJvg7Kt7WepAMsO4fESxG
7HGHo/5EPpgV+jvOIp8hRWpgLxbH4pWk5O0MSBee20fMKV3hWnGx5V5thqwBJL0VtU3qlanWeEc4
OUbIMOCUwn35PlwQNH9HVVBoWFr5qGEYaQYSIV5Ql2alg9hWjYvRpbDUgMZlB19K5h38gnCc3e89
hrrQB2qHJbYnK5rTIT70+qIx5AZlIMs4+FthLgtIsHXbEMVCPmivYvpMSuYGVeorVlAyZgnJGugQ
pzqgw52VwTJtPBDff+yEpmbNvlXBci5QPemrfq8+On5zllCKCML+YflzSAyi+6WNynaVXRv17qvW
8Sj1rcpbnuAQkGpV63jBub+3q6Js8aNmD+Nh7ilr/RROazxAdQJQ8RckimGO4rXXv4WbHNHR5cu0
5dJIT8NzqaQ1A9VoK6s6bIShdcfEcv3fK3FC++DiG7lwfQWcbATfiKfKI2zLm3DFzVuUZC0bCEbE
9Z4VD1ymELSE3ea5ILD9DJOj1JsLQPA2sysRaV6zwta3bXeYPxsP64Vn35VBsJPO8RhtaH/Y/3QY
p/YYxXiHf2eb1GIvpCaDo8ki5UenfQkZU1cn/PBJFXIbezJSpDdDdIsbh2Kj6g3rgiytJ/6fQjO7
J+VF+hzc3HkPv3mzH18cNE3z04y2IWDY2WPyXRio13/P+ul158R2Ykx8DX/7X5WHCBpiWLaYnuSA
C/06bm52paXwyX8RpitsUHA7oUxMZfiWNdQn2CshYj27ZXFE7jmYqLlBlHHWAMMhnqWbhJ5lq62B
EQvoF6Abp9SMJj0BOEysF+02+65WEL1k5f3HYmABRAEGCaawbwEgz4ppUjFxl8UC2s8JwkNP5XYg
uEMqpm0rI7tfDbUc09VhJMxm2kL3AXbsfDWHxWUnmWyUiL1RGzM7EAs42uaOL9XhqQNjIQ6ysL8u
EfCT1Wu1fdu23b0LB5/OPSFIkGSX45sXGJ0wQQGz3xfZBfDXuow0FrYKycWlr8zEO7qNPe8MGxYB
lUC3wCpsbQBSKTeX0F2JBPJaR3BifkXx0IrdQ4o65UBtt2icHYziJgbuS2u8un5KPrg1mYd7QlXt
uVVf/5kMaUlq4cEEdWuLx14WpAR0tI4ooiezM+NnZXNPqytH2T17fHNdOkL5VZD2lxx7rOnfoOcU
hcqc28VWMTPWQdo9h42DnQiBurB4Fmtlad8gEw2zggd4ZJKDFGSNqLjnidtqqfOGrsxLt+YHVI0y
2jEiyg4Y5O2Iyt304gTlxkIzOGcI1YbqruOX88DyZUDTkQszVARzk1sM1Z4HimZanKM4e1xSbwWK
mNILGQnrShl9+usYPj99SaEIw4qSiAvDfKHPrFZhpBIIePHpCe7F7bGH88hjGKSEvTdwRyi2QszV
+7wg0hGU5FDVzVP6VHUoNIcAB2upUIMHZXpu5074CvEvKBBrzI67iL5WJDyf4KIEL68sVw2E1P1s
AOfJF3t0uwoy1b+cgetHBug2MBur6DCNxIhtxAFCtCiPWNu1cIyFyKH349+Q518+kpXNCBeprjSO
VGIO+O76ZQUYZULMrYTQxogDybtAmSuKS53pf5Qh/WIkQx0STf6tOY04ppYNlfsLEPl03TtdTEDo
v/HM6xPU2Eyb3CD4oY992uy8Zdluw9d5abojOYpGYEsYqRJZstIEdtkGAvXKky4iXD9K5a8YnEAm
19JIpPd0a/r0LsRTZ5jE6d8VNnh/TWq2BuI9T1Vzx8kbX/sOE8ta3XS2etJMRFvYfZN4d9tlZqEc
n+QtvlVRuMqLkSh7/tD9splhAkdUMusN78kYg+Sd58HYiEY6+ljOBdrV5x6o3XizG4mXNJ+56CS/
YgC3MUZ+7ARGT6MOJIQjmVLM3yurkmaR39oVGXGwuEVore2hYh1BE6QvCNaqqopc9i/jOiU53bui
w1yLZlW90Y/WJp2ZcZSFGkSELahkWMA6c9Ti2Dhu1Xkma+3xTk9WadYNAKcb4j+d+MMcdqrDpPFF
6T5nDzxtFU8AUixJB6GYdatVs2fLYF1HfQLrOl89FSs1OVlGaNcOry86zvqEc4kw4LKCbkcQlDWy
kEL6Bv6pyyUc6lDjJfF5keYSO9Izfg9wjLgrLEWjggvbQH0XolQNrrWdbFr1j4FA7GB96HChciWE
/lNQudbucGZ7MmHrByVUFSTDQGtPq9QgXqEh0YWOwlL/lqZRjHSE4OD2U5QUOTqDD4jPCPp15vu6
4gh0PqRVrZBjx4yloAgIJ2T/KYeGjngR6P5NsNJGS2tA9keieuVC1NP5YOXgq44yu8A7XohCCXAa
f2WajTBuC+7ULiQ1m5Jbo4bfCDMUS2vi6OpmQaDNuX2wBH1T9XojS2LvHaT4Y0thlQM8vtK4oWJ7
++AfXx48Y5e+JNZlFbLQDTD4tJQIGIq84PJPdhei89Mua2iyYboNaoq7gi7LCQaW8Lt9GaWRRaxY
/ZCD1TXSQD4ddSx+kiUpuYwrL8TFQMPi/sTv71se0GPu0S9nBghWbzAcRMPgqwp/s1/wYJfSayaZ
/WBf2Vny4TCLaQWcrqRctcQSsI/ST/1/HP2SDaDrKWend7wZAxbvabw8TyuzD6bf8CS4Ok9A99/n
gXmeIii/2efiAF3Zx1ZApcXGZZB78su/l6xxkiYoIVrrDLk62YdekIiwuUzUv+zWf+/SEJ5FbCam
zs75nhV3Xxw6DXRK+IC6mBunWf5164p3kLwXe+7y2BXTqBSSoMHVl304z8SY+rO/7Cgi+F9wDAeM
9UP6V/AWDm6iV1jX+l59rEB7NCe0AVqicZLcNj54RUmj9aA7KvYvjLDIqmSaoKzg4zsO5c+HcxLa
DzxiCvC7Zv5CNj8CdA8V3diCiIt27TA7y34cO/hfYT1+Olgpsg/r3Pdsg6fKP/xtQUMzsghKldeB
gPUS41HfJC57VhwUb05W3fPh7VLa7GEFV8vT2tipSn7zcWGc6BX/qF4eZgE1yLV0k6lXd+bzhj3X
7KXZW44aMnkLS8tD5nOTSG4m5AJFasbsUBM552Wg3tL8D11uU+JeF8A+kYbEzBxuO2X3+2AKOO1a
buYYKFQdmO3V9KHvgSUz8oRg24IWyL2JcwCjmlgzfafzhmfoDUDn/a87Bf00L/3TK4y3oismECCC
jy31zmUmJsDIl9+1Z5vWgX2Mabxl2py0ZRnyeElUxFD8MpVo0+ahJFU13G0PYvQ31aG9LAfRAbdH
TvuXWCIO4g+z4rb3kndka9szPC7kDU4WENFKJS9LcSVxO+xsfd2vL3SEPSHqEuQLInScSEzQZaAt
t4z0uX3LBiqiPI55pk+4dRWKi22EhRnyL/8GOb+v1/ZipGeolgJhzo3KR/8DeMD+nt3Ka08WpGmT
ZDplqiH02lXUQ67ZVwTGBswLOyHa7KimtGRbgckPIbYdnFYoXBxGgirU7Vib+J7LHDgfi8hn8mlC
RK/l70T5kH16UysWmsbuU/ExQMwjpYShx264e5y7kEOXxk0PYJgFHciuNFJCuMdqYiwl8Q+e3cwX
jAImcZ+a9IHfq/7i
`protect end_protected
