-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rr+ijfZ8bxKEyoJ2nRdy2iGbERQbndcy77WEpqLwjRin4I/dfDApOoRjG0Mi87+nbLxxK3JRCnkB
p/IlyJW/4tXd13CMF1g1S2tal0FyOrWO4lqzCskRmFGbdpAntFdLEA2s8xvWMI60qVWbEIWYCXxg
3tVV6VWp922se4Bc6zeYLyeDQ/tYsN1AyuCpLWjI4eXnrVXlLRyALh6NTE8gZ3rj1FkFwwaqiI1o
exFtvVYJfQY+geW7LUKW8xU9++WkE2nJNEoAcEf5RDZpQLYbBkDje41x4uhwemMzctaEFitNj/Gt
IqHuhrpWNbTUXJYuu0sQbpmuLquyFIwvh1RNdQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
NBO+l/04NvyHzzczK0e1ziGdqPdS4dzj1DzYqN3yAPyl6YWp19z2iDWD1xq/4g0CRa0nbjoqP8C9
x0TsCDc9rI3Q8dcCXE6hWvNjYIrzSAbirqdvJvu7hXO/LG4FIV9h0UeiBmBPWEI/wLQyGdLdFo95
km1Q4lhV4iTpC+vdo5VYN0FCGxpYdfbavv2dxujgqJ40QrcrIoEOvVvvaLbZDT9lu7Iv0HHWZkEt
BcMN8fJrfAmzYC8Pjc+HWO4O4gkM40vUMXAkSkqXB79rKLDCDxLFAdRIJdj488gyxO2zekSVgIqZ
bIpPCS3JVNZwWTP10RUm1N6sjLcJ+uhP3u6xa+SaOgCgDOdyKp09JPw71OQqzdfh/6nLhhe7rvL1
Dc05k5DGGDQHcrP7xxtW5+DvYKEHc3KVd1H5YIzB4t27F9FUZZM+KfBJssxxu+N0no2DRRDLqhkE
MTnRPoykj6mMaJsf10Ysp+yU76Py3SzRUV4erbiFB16YDMGzGAienCdzAb2Be83E9QKxkL67Htzt
F6RPPZOJTu4kAEw4h0R/2l7NzWzL1gC73uvlxEkGXx24GZGKlfCUkEK0iEgnSqy6V7zkEu5y/rwc
xpbmy2p0h8tvas2IgpUXnr9SYy0dfGEiWV7S2L1azp+FEjlHvK5y5m/7GrPTBXIF4iMmRI7wAVDv
UtFwhrN9XX+QKmqkB7ftKMFF0UN+4ITNwBGtoQx198k/tpej6G0wlNUbNS3SsqVy4iL5yB3CCtho
jlLJjQqLf39AVelcP/HEEUsP8cn7XsFw9KEgfK+5mSawFTU3urPV79pRvlAUZ/+Vh8AvwRwYEjYx
UzX4oD1jD7GR9lB6Q+qGKU94YfMiZE4Gf952y784HFziwUROUxme9AlxoJwxLcaJnJwm4CsO8pWv
/1NvLBFBUktoHXDuFwzoga9ixJxeeaL/Exv9vi+NIPPzsQ85xlz52s7zwbN3Vmbpvfg/QtnXE1r6
hIBwO51XwEcaLBHq6GyvPeS/HWat6SDAu38bBFY42+N5vkX9RcxKxS9Ylne5XmklnhHaA4/wpJDT
d1SzSmFG7CcE8j/oBWmAbC2HUl0+z4DS/UkICQSOGaAaGpWVH8T/UK0Q5Rk2zBiIngEKOBBgBmLY
5OLeecNzMQgJTR6EAXtxMB1llwt6Oa/4BfC1w8R8Z9RFmfxGE/kDdM9TVCnR9tCTsDZ/VUfvIF4i
lZy8+5At9yWhv58BboOS/rqBSRumWFmcD+8VXUv85RUComEjjwWd59RYgLXqnF/rNUPWxqcO2Tvq
TeJ62I6CAoTxlWunTAkWw1dJKXhQLuiK6cMWIsVPJB29nWIPm0DMqZrnq7waSruo42CNXvbiaYBn
RPyhUP1SApgtkjDLGXSSccRVndHTmhOVqt0yzF3EdKPrleJq39jo9QL23OnqO1sGYpC2AYF/9SF4
+E6lzT0+GqOGezXxrioWv1w5zMuFWsmEFFBaNkVfYwSLhrmmMTx1/v1GnPbUflHNvGbTI6JjL1iH
I6PCgacn4HVVl7LjNwji9B7z+PvDzxtnmXC5b5etZeNQd35QRwzuNGISCar3C8c6/C9ltju1YvjQ
bL6YcS/LHnd70w6gwDEd5yUvise573iWsHKrkSKigs8ST9RXC7DR/0GQhEQL/R7S4eYFnP3Fc0ba
BAxqrtiaJFAjqJ3rvGSmMbOpvtRMGYjebQAjhdKAP4nH2/rebsIeGMwqr78kg+DkaZIt7ZanSYm1
4Oys4obEWCPTcHYCn4oq148rcBwtAMpdQvqZa0g0Wi8p35fLs7RYj7326oZ8zOWY4ZM0+yN/MlE+
+7y/nh7gBkoi/sR3VUVScoBZ/pOX54OIkGUzaKyP7CCeEYdx/9ucsRv5diIWmWRewMNoKF3su9Nu
bk6sBlqwBnF/hC+Vtw9NbRCZvouflpm4Fz/UcdAffbJmbiNa4EGKFbuE7/Psojb0y2ApmwpqkADI
zVmCfT6Xqd2vt0bbBeBQyj9Os1HY4+2TUOP2fZUaoj4AryDuPCS51PySBPn0GB+sm5ahKLvnZOQ6
GWW2Cs70FsG3LlBr94Uh2CB43OxnjxFwjtNowYhAcu5JSyLpEKSHd8ZCjh2PQIyUU1C69HZOwWVO
RE6pltoNoZTai0fJP2N99ICKmrKQZ3iEw9+FyTiF/lLh3YSHOKmP9UpwAQUvaqJGoTgCBJ6CMRf7
Mu9/MrRI3AVho9QL0YvfBa3J+MffbkP442+3LJubqvil+MH6GuQBIYnUKz8Vq+qqiSuVUXYwIxRV
4lrSWHQhaGng3DJkh/FPoTEkdIl8L6PGcEIs3h7us+ecyuVU8BylkBQr12JBVoRrUbKAzG7Sh5zC
Gt/OHCts2MiGE4I0CRnMAp5NIgu4FjwvReh6FEMAlABqbPwY0BcVoJRqW8gpA4VkQ2o7s+DiElpf
CW9/tzTwDvLy9d4r0WXQeVIrQKkx39P2I47mmTcPqPzj5dthYF7+Thj6lsjW+YvXOLbBkIYAKJ4z
zWb4vsDUbz58ds1vmiNAWOWHgIl2AB4b6WhQ5RHTzOvUIDuS5w/IFeiIuANIIWQPmkBONLAN8PH5
OdAhLbTX0eS7pQEUJhaowO6nn/kfUiqT3mmID6jlJcWqgpmyp9COmWXMJ9SPM1U8iDhLPw7y6GPK
+EeAmgwN0kiiuJm4pT8RUsQwdRB27GuShtzbRfvqthdGKRuKkZCN6m52PW4Cxeh4K/C3C1SDYZt0
xtmxfXMbK/urErP0/GbICAX0c9wM53K3YoobE+N2BrhlmDr2O0hiGimkjq/NmzKN3T5vbgxz7zSy
Pvkmb28wrTn0H7M1opWigdGmNcwawKgGyPFX3W8EUDkdQ10pOBitme6ZRB7dtHzQBVhAvdrI9spe
fWojdfc2TePp8bRyAk52Q68e3f7aHeXvz0jSXBmjphwZPDyUN1LSv6DEJZVU4Lhp1Zh3wdscADXW
kKQCqTArYmzlz6K6/qN4lds5EmZK1RHY0T2x4scbdlxtHmNXBZYM326HiqQHS5NzBkCYllzql8lc
EDMWDQLeBA4e8UA7xf9fM9lW16mg2sFdAj/4vKkqRJ3x39nkCFQ3dJL9WWW9zXtGRx8JExGhK27h
82AvnZ9F7o+RF4dQVww1ifYKe8c56LpE3EydQK8xub1n9Wjy7+TiuZ1Za7+DbQkdUrmCXzYW24rR
L50A2tHrWHDTKsGUJyfIg2+rgOzcfP0dx9kpHuvbs7MhiloTfKpIrD4PQYtJsHq87kKVA2FWJZIx
J2mrhwC81WWELxjoBfqZN4uz+vvEqf66PuJ2S7P2ov3yMMiZFTlTAhXNiynmNU3JsrdkalsyN14V
DX/TlAB2IVR+TOKDRd1A6zDq/1ssFAdDUgTZFjzHVhKea3XVSWvza4q954Op8dY8o058CsCtYSe4
ZhomL1TPVD8W+a9ssWj5xWSZSXA1aybpUQO9QbkyF7N/OCqg1Ii1oiK8c8UsBHg+Qlz2uUlc2IHZ
i2iQoj2DNcw9PiHluPEizUtSRXaP1oQRuOiMv5UbN3MDmN2rW1DvkMAtQQJ9ePktgEhKe5Xtbzvp
Lu8MNv9tKUMvaZpy67CMmcasXOouPcM+kyE74GFx+wksiSZVjTLBdbXPUD6BQw3bORXp1T2B/ME2
zDHOg4g0WDstTypbskAxNSPDmIk/cFXMJV3fmTXOvIwsG3wr8++2n0BbcdDKJU9Q+/gGISJTqs/t
GFipgybNT3GdBD/Tfj7Nk+VCbqxG3Dw4jKKbrSMTsQCJdwSlNDFMlPIBVtNlhloNJBxR+KoHS1+6
SZDyQ2rayEO0tsM0All8i68qB9hWJc78NZO6FddBkF6A7Nn6NQoW2Er8VeM4nS0zfARBy+e4p4OJ
1PQDiaN3As7VpBW6m/pxHXtjeICb/ZSehr3e08kKlonPXC9t257r81C+tbVJeZbD/c6ze2vclcO7
1IMyrHE7a7eYb1NZgXUy9+RC/UUTKPaVcjHSPvY46ME37oGNksDvVxVWBhc3TaAsjZdJQPJZ7MFP
BF1ozG/f9iiKQDRXuKSsMPggSywrT7mVTMRAUjlO20qngBEfVZzLvSK1ItBU4MbWE5owCyjlpIus
lk2Q/27FneMRmWXqqIYs+tS0GbPb04S4oxjcqiuQL7Z+cls90C77/xQHUyJWJ/qFqhf0OQmznKjt
KuBxRgeZvp3YzRMquPd/cwX/7dUDsB6MnQ25BujU5AUQNZwethaCCxY41t4aylIxnzEUUqxqHjMA
NFI/yueSIdzxQag9xE9Ita88/xcbVHhAjT0WuVZNr4XUIzi4r0iNceZSjHSXJkj4rOycYn/og/wa
RDi4yMiEBhlY91WBeY2rYMtZHU65Ip1+OLkVFPKyjnCubLKhgaRrzUH+8+ZQSu90ZFTnFsnN3BmD
7+QuH8RkL4vwN+wr6xvjSdiKDarHf0fcOvWRO7kDB96ohg0IUIdErrKKmiCgZhlJYkE0TNJsaIb3
/pIZyVXtiVSqRIC6iYlmP9VMLgb7XnmvDRTmMCy94xE0LG8UZJFkU+rnMgXJuEUC16o89pXceOjW
bAT4sBtkSLtSmU2ChmR5hR0RxktAX7B8tPqiNqqlQT4cRp0Y4xT38Bv/gWG3NSw2x9eRcXU3/pED
F+q9guIbUJK9T9LZa9A5l39S+vlf/0Ga0d5RSspB9+jxzAxhfwlXY8Xbsz2sIKK7DLJ4ofFR3w2Z
xN3wOFCv2QyzsEHmaCR4m11I4gvqeG8QL7MigF4UjzynUu1RWX5KF9ZWWM45JKLl3fqPPf5SBmHi
Y8vZtAAfD243EUwOP2gWuRxBorOV4Dr7yH5ejkus29loDTreaEeo+elZR/3lJn10zsYC4wDmZjnD
CgCX1Kr6fvm3URMyfq3ajHphVJxGN8IRwhlqtISSgh+6ipcGs3/f7H7pnrAgxWqchHGXoKWOsync
riP0QZFsQ3q6xTG1n86xkbkWfzkuxsyLBSILmBNPi/BhaWXUBtXcKGhmim/7VeWN+GE4Mvnfs+Xu
KAGYBDXYMm1049YEYJhhYi2GSGpIgO6FtW+Qwu1bLqKvdcGgizv7s8VpyITXlFH+2oU8cGilJYGd
SIYuar/bbybEY3TdvmpdgGtvN9eGR4P4E72ArhBmclEtQasmjfL3eH0x78mCFVRA95SHlItSboro
DDelaFvN/rugEyqeXKRR69qmJmP4KlTDagujaA/AC5RcogbMs84vu7GFblWlRwtDCYqWhlJSUY6k
fez32uvXvEysK3WzfAiWGtrbb1rMTAdK96/DvZgUqO2EeICnOEIZNV1MrY/J+yKyPMOUG/1OBgjr
hvopBwTbk1SDaP3o+e21AHVMzFsIW93n5ajs3wcHToHx5nuJIay2/+NKb+D8iA/CwzF6k+NV1lC0
mNpfpAEBHyyQDLct5NRZSLZAZencMBAAbCTynfk3ecZshQAW8ScehEYxpcgHxiOi7/TSNZ9VmyUV
CdOKo0b3drRoiNzdAu+t/cOkab7djQ4HMBRHWYtHwYUIX49DryjQlX9k8Dwa4SW8psnDQ4/ohYYj
U+MhWem4jSdlREOJIqn+hbhxpopgPsW3kANHJq+DjnQ8NFeo5e/pDH4jJh2Kad5FHcidxmLgbi2G
RvNXIV/mdBqRaxV3WgimmJH6wqTdIDRjBq2cgdZBXdKWTJ9dLJWd8wF5WgoupqOe8qMTzE5uTFO4
6w4D21Vrq4kkZSfPuH4S/Ok2HfNZzgbGXU9pHahNsfRST4bSZBSO6sBB2yA+QY3mOu7rKO/pc3X7
n7PC5rSwCKKa3GW7zYzzF554aX14PReX3z5gejCqswvrCUvF0BaVeDOR3DpojNOYlhtYu99LGoUJ
eNbKS43HebkL/73G7PPzG5t3J1hwetxw8Rgh5FkIJgLfLGUIXQQUtYSOMrep+VTTUti+UQpkb/hV
MjA3d72ZHRa2iaRpGh+/cEALq/gSbIsOfroKCDQcajadKVfZMQi1Iu075pSIVIgyJoQQVUWhC72c
eLHXrRI0lwDcsHzJqXFnq34MkjL6wD5UmQ2gna7xP8R9Wx88ExdJVu+ASautNZQmsLaWiBOZiiOb
RoELhlegQBD4HdIpjPvDzSBJZ/cSqzimy+JdkdAtQd+2MOGjsAemWKmFpWRlGwOPLeR/P/rgKQ+R
8wydwNfeWFylR7gsRRzK3nE4FnmehMZuvezRHFMxRWXuWuCWrxZqi9pxcMC6oBOn+Ss/2fFPa9kc
Il2IW+qDrO8oE4u+R+Xb7I4H74HbKZ7gwraXkjp0gMiHfMbvRnPrKOzXA7AyXf0Rr7+kzB8/3olr
BDkr24HPyVYu/nt2OnbfJB3o8skiU2oZI1p+cUuRjF2c26Yjxm3bERXQMLXzvCKca0UCgDp0u2mB
PCsJ+8Oy7Obk9zL1erUg26A50msr1exKLf1TdXCVJ9vHgBZmWcmxo03PC6UtrwPMfAp/VdjbP66F
+v2HoTi7G0gK8KWeHBfIf+CX6GgF7akC8eZLCpBn7NBPz26ocNA0Qsu2h4g+X4ikwleXVwBv2AIi
H2LQBa11ESNt06ZphedVUwjqS3DA1EMKfFF2nI4au7YDugqCPeR+NJHWIExijDsYybGH3O3C9e0j
J5T/JdDVmOwFs3WJfHg/yntHpCzMJXZV+WR+m9VGN+0zznZ4c1YvBK8SfT9ZQjf8bC5UB0eHv+hQ
6Pcsn/b25Ak+lwkzlTDNa6oxbsytcx39c110nDrQYgUqMG5IrTCPgiLSvzoDGUkmPqZ/VcUuSsnz
6SkRKCdbnG7RB1Gzss90g3PWjgDGvQmH53tXoWZIb+1EKbFWm8OPO4Z0POY2Rq2uNxDlme3RFviC
UVhIADOP9xX0/sgXxx8/wcd+ztT3TrTF4M6xiFD8986T2kLuZSJ3VSct94JBv1RqAy2P9mnoa/x1
jpDLtAZjtxikvIXYpXVPxWxwXM77WrDpOF/0N9lEhx8H9diiW+RpL7BiR2Xm/MywJhvYWioxLx+k
P1oVNKjQU9KMsI1Rev0gqzbIpyH/PRBU1DUg0TWrYopiQbnFF06WQdUO7RBs3jOqUk+yTcmeEe/h
DaTH+7IB2JcV2FEHYuGvYMkRN67dVf0VltW8VQRbyclXTsQIb/Imsfi3VNt29iwtwEbZs+MP2wGj
NtkL/hGxb5NN6JhR2mFzvPCtnHoT7uV9HsnWekgVN9KVpERgBJQqm56WJb3EJoDeSV+Uf1F//WKf
DItv6vREiD1ywaYF3sDTSdiw1/omXnuz6nYlGadPni9cFlMOG5m88nB01wDHnsk5yXyDQ4RTXdyh
RYPRXNYVYTpP7VhvoNhsVvi0/ABBR9iNbG3Ih9v3uYaAQ/tDJut9rFA2VYWiK6IuTMCfOGQvcXHv
4cQZvWt1KS5ZyJ8etiO0oqtCJX+qlkcRNqazM+j28v8AXTvvsXLYeRVVzotlg99xaspKFF39yAOk
z5YBaaPGoSsgw7pjbs6iQ5+s9j/430cVmvkTKiDwN1Ymsb7mVecwt/U04hnBiQOMeWPikQx2Br0/
tFLmEbgjULux6UWHLqtWovXxQLaHdxveFIFxc1P2PvdDyrcnvxK4IywH1g9LTsjdXkBT++ZI5Ctq
DIFE52DtVRC/5sb3SpfqqN0YMEuWGIf1LWPAlxbW0Yy/inJjuRt+BLhlerTj0AY7S90jjvGVN6+6
og4Z7pHfDP77yGgriPeadAObN5HBrHcwE9BxE2soIgysYyhHTiyS54k8Z55MDm2Bj0wimRd2OwZb
mUwRrT1isV+lIACOlnMG2fHw06ao3Fju4KS4puN6EPJqHoVD6bFlbU7kKQkBmCjddM+sK9OBVOAt
9Q+Xi2m0MYOyaufqRZFZKHL1RXjn8fP5PYIhyyjZv/Y3P6QVMkzhktxDCL3KeXjmdk/SUhUpkk7X
edvtve3h8Oc+Yi6b1IQX5R63U7w1tcJHHXak32jRZsUwD2ZTPx2PxKtExVzG7VOH5/D9vRoQOVhR
MJECkF92CqT7a+2Shta9Iev/jGXS/DQrEoXJiRTtIkqyftkVBsJAXDf0bPJsk8WXz6xhM0HDESZP
fzgYDileAh6BkrNVgIrV0/uEYkUjEC9Z+1f62haM2avIV9jYhT4ruQ/IdrdMYm+ZbgpYiyWogk6j
JrG9p04LO5x/+cuh4bPrGMlaKxQM6388zhCS9tNUWJOPbI5zshooLlCIaFqqio9Aan9mrzodlxdE
U5e56e5L8bRD9rR/O+XhW9lrTjRKNbSkPw/3uk+yOivaI6ATPlzXC4rW1Z3s8wApYuH4C9KpWb+2
vc8Rn9CMek2qjYltLSJM4pof8BGw8T1HamIXEpKfQBybCiWZ0+3L/p+44CPf3AjExMgpnd2fzhxw
6KtCIlxf0KbYvqtLW6eb2xA9z8HYj9LA6ZWGg62eabyJdMpt4DHMva9IX3uDPIIiPwkW+KAwaKNr
eZ7MD6N/vs1C/kXoGZ972E5a4jx2pgbMwLB+tcMhfJCXPm/ILJo74KEpI4rUQBVpgizh7NN1puIb
81oBkH7H0er7jQF6CzjFI5AB1gTafS4qdtakdSdZr2HAOkhKxeiJdm/uJmhtFKLjRZ5+cBPtPpcC
waJCNjpzqIwn9lBaCa+2moUqIr2kyHCLutjPYvJhazK1icY406ihsReI5CThf6/uGlVv/+3otWfw
IJ67tX9/vh2tmkBPhonOo/71GCQYzQz5yCw8mtsHCtSz0Cq/5xK/0KDgmm6i36cifDxctaBk9i4q
lJ0z7fX5LdbFerBO2UGfOi4HtvWmOjW0nl9KrVZepiaWxbM5alfAzM05KCrK4w3zuWYVNGOZTq7x
I7CeaYqbGnHW53XA52I3j+kpyeAkeEFBFi1E/Yw2kMIyR8woYZ4HVWfc/7Kwte+mF8UBKiu4h+JT
SIA9VpYVuQ5DpS4u0diBRimNctjVReoAkvlJl4U4qizylsDPEJ3nMY9nbWu9rl/rvErP9C4oy9F4
C4sTux/76ieRofka6pM8tJNUEBJH5Pncusnw1AupmhQGRk7p7hals7QQMM4+qFoKOrBgWIiHmV7b
77xpQOVJQIuKxMn1y93uOsbN+5Dxi5AoFz/pRpPcTxgaBsHXB1gGwUDh+l8BkJJF7wP1GuUpfl1j
Q2BjH5ctAtuIYs0qCjXjmNTPODCayTUWxYZTi/DgRDsTqFGyagB8d3hoaIAdDTyMoztXyPf2EKNM
X79+wURvZNiX55txKFiVmmVt/0iBNCutwL9uk9Ijyq4BBFWB65iXyCkcYio8tsFFwp721MOgNMsI
vHwTcKMY8SPMzZwvk+QAzbfGy8dACutiWxJvNSHvtvacMKcxHqOdMF1Fk+dS4X+ApCuN7rSurVxr
DOg3CxQzu7yC7yTYCpzMleKs2JxNAfmI+bR9j7hITZN+VvW55utlOVbSwfVcNwJhneFRXZcDUyCD
DjQOdwjzD/cLyawFDdmxdERj8w2dxlVJ8ebjJyhEqZn60ieX1Mon12SHlB+GDvXNvhU24Z4oTHti
CV5IFD5aBhdaVAfjS2xPBTmRv398AavNvp80vUFRAz0xd7kUtfU8BL9ZaPFaIg2R0uUcfwv4xT0T
gjrsGeDthhcoiP8ZAPhdYbqz25Lg8XYqg0VghRJWCzDLvzRMwSj+F0XohGKbEWXcO5uizrp8UK9i
CZdYKq81fTawo8a9H8a86iYnHX6ufRNO2UoYPP4go1/9FyJBss1MdbKU7fVSqn9jSMwE/PPeyA2E
0aX+HxRhD8ZlKDNxo7gDtwtIL7KRLo/JIBaauICnfRR+s8/Gw6rhwZEdy4fpH7L2Glk0+4+d5A5p
ZnneAVxr460ehvDFD8O6zX3N/k6Fk22hmy7mfjy9Y52ZXENGHtpiNU/F8lKhGgwTT1LZ97AMTtJy
AjEt3gDKD0Xsc769XJJJsyRGqgxT9EdjB+LwZ38zN6TnYGlurC/SgW1svrpFWGwoY99v67TKJGU+
LXMzfOx1XeqMqZ7SPucQxkwI6+t2EX9JVLAZlmHEpbR6ALqnHvvDHFvbkRPlRPpq3A/3mF7jBrkf
GLv7kZygKNWWAb0Dj/RpMQup9SbVFrfnMn5dXbEecxMz4NUpWCVTJQxV+gTAb5BZ4Qeu2wK634/z
3csFpm984vUMpTdcxXDoeAV2ZQL4yqmXeVMxhLH9DFDJq2yu5jGieILjylOr2WCU9//mIZM0Aadq
psPl5VZ5fIcR/tE7cJ6jqA9NPIdgsYFNIbmci8iR4mjBBa6OWtciDYpXRGKuPKuPgAhjsGAv9kAo
FwnUkObEdsuWpg+CF/vS2Na/jySC0zm4hGno2Kxa84eJRLYPYp2vonByYm6JO2EsnAUdprrVzbGO
F2A3g/aMmp28sqtX0zj4cN4DWJ++Ww9xld05MLuoVhElvKb9BEhqTtYwrFWyeG1WywZ5VQAeuTCu
kdekkg/NQ8qU81d0FscmxsbO7CxMbJhBOoFsMgiQGrNGzq0J7pHhIOvPIne97UbpDXoFhqjnozv4
Tg34rLs1L9zpFOIyE8JDtpItSLPy0ZNLxTj4EvPe0ZhCl5kqCUdSVRZkls1AiApVHGl8YQNVAPcv
GWA6kM+CsZDTNmbH8hONEBqSUAOeivx4oZ8yzmZ3i30mncBPxMKqxoxAc99i3QZJpRU89hafmmHM
U1G1etxmIqwxiKn+RPdmhbUhSIu3mqKwx2s6R2NeoHk0JVA2hKktTBNM3KWZvcaRmCqONVYFCKHp
GPvA8ya4NlJKGleZwAEu/m3Ub+Z5saA86BmMgOEJmg4gumv5gHGx1G/fHdvvtF9RhDytbSwIFY1/
tk/hxisRfZZBE3gVrxqbofYl/JfC+Ut92u1/klFaK55XOhT6Ij2cu4AYKkM1depNdKe4zu6A9aSW
2x666bFlYeHRXJFWQbXS5+kkCBSG8ihGCSC+inZEq1e6WcuofdRxTPlUnCfvBK/8hChTWhIonhEW
`protect end_protected
