��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_�>/��zTg��P��Y�@��+����t����m"�Q�e���VW=I��K�']��GBI��|vz�ٸh��?8�2փ�%+.Ht���P��D�C1�˟L�<z��0,�u�UIj?��P�����Z��WY��!���݅혫��:��P���G���a�K�P��D�"0�r�,g��jߥ�.1Y���迅A澅��"��ث��<�X�Q�M>9m���F�kd�1���ά�~/��1�Y;[#K�G�J'����`˩���@\1�r�=Kd���Ȋ���q2:KZ�Fu��i/��%��;�3�����f�D�hw'�ˈxl�t�=��e��H�"�c���L,.�G-H/<��)��'��"�u��wȤ�����&�;��Sb�A԰��5(P��f���TW;3m�ƭ�(F���|�\j��f��$GN�%�Y�td�_���гHN�ҕ?�4��/�T��+5|�G�g�ʾ�W#G8Z����|���䷂Ea֟VY�͎��(�؁)�[HnK�е���iR���A��I�ZPM�z6��2��R�H�c�@�J�&��h-�������0����H����.�oH<�yS�T3,*,�ndȂ0���XYOW ��u�����q�����>�E��������A����'�{�Nݗ��_A�$"_���J#bD���U�ʮ�a�8������ L1"J���s�����ǋQ���8m���%���̄�q�r�C�:Ϧ�;1��-�Ŷ����K�'���<2����^>�p'C�G95�4��Zߵ%�XUDE�@���E�����lߖUW���o��7Ҿ_d�>����J��� ip��/0�Dxu�[%R�Nu��ȇ�mM9U�T�I�w58�4���J ??���H��o���1{V�h��_�1Y#���XYv��Pp�{���DĞ�A�� ct�Nڅf���\�9�BrNt�P+xne����DT���6�V���UӑqH-w
bҪ4�G���i� �t�q |1���U.��&�CHRun�J�C��zq_��Yb�{1���WSt�����>g�e�F_a�6�����I?�z/!��d#&�c�t_��@kc&[ɰ���tW��)�
��V�N��F�����}�i�=���J��ڤ��s,�����~�뵪�AOYHԇ�
r�!xk�T���M�6������a�M�ѭ��>A
�!�-Х�@U�Y�+Jj��w�</3�!�Ucyͩ�+��k�q�z�����itw�nn��\{�G�j~�����(�7�8���+��+��Gp������"=ky󕘏�e*{Q7^�)��,���|{7�E�Dh� ��Q��'����|*��QlI ��t�st���r��Js�<�q�v%<���A��j�2�w��D�p]&��r�v���Ib]�`Tjض۰���o���(ē�
ܟ��w$14u�8�x#�Țn�[���� ���~��ۊ�rI?=����i��@p��<݈7oU�����d�������$~��JacXJ߹�0���K6H(o9�k�Q�l�`���'��n_܄b��7�4^�فey����u@u���[�a�����)���nY,5J��y��厶=��Cz�O���ӝ�uf:���ڈ��D
N�̳��Zi��c�Pq���	�c���R�Z�;�.Mv�C�d���̼+�ꬃJ�	���o�ȁ�����)����:�7��,����X�_E3B�7��"X�4�+��ܜ8‚��BCja��n��G���	����x7���կ�0&g\�S�b�U0�z���;a:v�x�z����g_�o�yb�~���ֺ��o?}��`���MKk�	�������kЂ�)Fa��YT��w�|����z�ؼf�j�B+3�P#X}S�.V]z5�tl����9Ep"�]ſ<��ϫ�����=�Uw��W<������iȇ�`K����=J��r�1y�a��h�e�>#Eڳ����T� ˳�]ܿ���Go���/�(����u$�ظ��ʶ'!k	�C� �����	I����N��6��tv�=�:��V����,�)�I^!�v�����81A�}EG�i�5���U
r�7��V�=Q��`8��@@��+Y\�Y�N�G�c~�	6� �1:2�2e����ظh%F4�HC߾�Ӑ�����.hV�&�*��Z���_-6���+B�˕�P�R=���v�qH�~AΌ�*��2�#G�L���`m��J���9:�Z�
��w�8p&d2�m`z��^UXH}��g59R��+�('�а�{�@:�a|�R��h}�.���G��������ffK��Q�(�2���`Ec��,����M8<Cc� M/��`�8�{��?SU���IT�0� :|1�@S�%��m�
+
	���󏟶�ݑ���3L�Zw9���W�[N%f��D�����O.,@NXj��aÐ� R�wV�J��k�_�i>0H�B��%~YWc)����q�r�-�i����Q�T�8Hg�j����� ua���LS���������s�z<����7���W���F��>̧N��龬0Cp�t���M���-]�}GL�Ƽ�^@�/{�h3��ӟ�ϥ���Ԩ�+_3�0�G��,����{k�z�K��5���PG�p�(&��s1k�^�u����jً฿�>m��b2����(�|�4��Ȫ�h� sS6Ȯ!���IR[� `?ȑ]K�P�q��D��
�p{�XqAG��d�;�ŒC��D�/-�"[ ._�i6y���Ĉ$4"񫘻��-�Z��x�o�~ƀf��S�ܹ�"�I�ޒ�8����x�DȰH�)\o*���X�Ň�[/��^�eR��pW��N�2hk�+�0�s�3����wj�J��yY��n�<���W��]�+Ǧ��
E.͏��i�7��:�jX��9��3�ќ��96˿x�c��:�r���S&V�>�=�j�P��͛�����FP|�|�$�|��<9X)<�u ��FI����*E}w�Di���)��=��X�HO�c���*�v����nhX��t��N�;ݏs���'$�����.d���
&�
�n	Д٫�\)�xR�&��K
��ry�T|@ՠN�'��-�y����g�����>������tO�2}���^��/K�	.R�r����r���?�`�|k�̏#g[��'H��A�R_Ot������2E�Vۂ���*���+�^#L��>Rn�8g���%����2��$RE�Gu��Ń�5P �1o}��B�W�}�>K�TG�(�jg�!����T����c�/�r��'�>l=a��S���=��qs���ي-�w�\�Mz{��6<�7�b:*��<��|a�H;���p(j�W��ϥ�N�tt�x	�����ƶ@�8��#���/���(��赶����@M�]�W��8j���2�J�?b�9|��/��q�N&!q�T�!�a
5�\ӧ\|Q�����)F�'͗�%���Ӱ��)���䨏֬c����
�#di��l����[�0Xp�����Ir��S���Y���KsZY�����@cv1PZ��]�����(�?��1��� �`V�҇m*�69�ݵ��c�R���(�;���BpY��h�w-���m��w]��~�x���i��@{yY'�C){�Ì��������� �L�d	?��)5�x�P��_
p�J#O[~������w4�׋eX���;��!]L���|��lh]j>�����]lۇ��3�(��w�����a](���9;��.3���ݷ�C�P��Tw���2T�-o�
3�h�X���=I�%��'�j����U-��y$#R���˸�O*����q������<���7��өۺBU~dW�e��<Qa�,&b�s#XsV��-Q
%w(��nxH�}���qug2���ﻯ(���+�n�(w��$_3�w�:i�=��6�w��j�VQu�+:�擉���5�{�,R�M��>�|�D���Qk��0��b>xT�����8�W��������n{�3��ַ׊Sc�Ȝ;zђ�B+��)~n�a�H<��nX�n,Đ�0�J&�7믵��(<3/ ƽ����z��e�V�-n�����FT�����V��5�ʮ ��֋��j�a��2hQda Q�;���1V�@�S�7,�x�0�D��F��A�]��̊�52��}B;ĻH���Pu��RՎ����k_���:��������xe3]Y�.�>�5�8p���{�9��+T]fL�
�3&'t�d#cm�x��c��C��t2x���Z�G(V�^�G�+�GZ�2��6�h��൧a���xl>),56c$cX��2���>�:���S߽P�BȐI��ͻjV��[+��To����-�5�aE�� nM��8L�߿�E/!�eC��nT#�eI9=�P��|v���ߊu=ͯj׎��l���*���TŤ^���	0����>�� �!��˘�*�Re�f��e�BU���6�Y{���Z5�^ �)��T�����5~\�6���̢�@7z�:�n�3�[x��	�t��ju��r��(�κU%a��T:�
��؁q����������7�7�7�1 �S�^_�K�EF�Hހ�4�`�j
�B�%}���;���6�,�K��z��p	��=����gЏ��n���ޔ�x;~�+�M�m�R���Ji��@�]�Iz����ű_�􈧴ԣ�a/��Hc�bX��c��'#x��2��ՏL;r���%>�j���m��I	���tͮGH�a	| k0uG�a�O����5x�I!�������_d5�r�	Y}�^�Ga�HoD����K����J$�?A��$t]c[��Z��f�h
S��]�,�������q�T|ݍ|�K�=s7U��&^�S9ンf���y	��W�8Md��7�h~7!�6�/:��~:�z;��rg���b���Po)o3�|*��Жխ�U��T�l��0UڝTYy��`���m?P�u4-����I�\�� u1ޏ���Y���1�Ü��+ة��Wىd�#�/��vےb+��ĝ��C��ZK�A_����+���_N�)�P�-�	����q?~�/��D� ��+#r�g���;�ؿuH���h:|>.8�:2�����朮�:��t�_��@)i3)|Ȕ�1�Y�T�-Rt�/��T:��A�pus��k
E�WLP�=�ݰЫ��>�9~'�w��b�"zD����U4�'\��k�v��w�s������Ӎj:,��U�-�tsr��7l@yu��$�:���핕���]S���6A0!9��K7��(�2�E�Q��+��b� �ğ�� �|��F��hx/+�mu�ȟ�{�n�as;)�EH�̳��%��gտ	�F���;��"�Y?�b�Z���)������q�٪���{�8=�%^��g�C
굑d�(wDߑgT�ݳ��M��G�0-���}�I54��S~ ��dyX�g_Ez��m��q%w�+q�b�	��[Ms�	�?}���ӔG>���G��#���ê��R�Fu�����=�kS��|;��VW��Ƣ���3�lA�8^��b���b;@�^ZnI�Cۖ�H�|z����}��[��S�?���V��yh�(ű Mk)@�c���@�3�&��
N��p�V:Q�sa#�a�\��XO�I��?�h�:@aA<u=�ԇ@�\[���d���%pR�q^�N�^jf�rV2�A�î'����$����_�6;�e�_��B�`����sGRupq~J�`Z���4�$� �U�Ȭ��p�阴ysl挝���[*e h�^2�� {KCƀ6 Eȋ:�h�ؽ1�}��T�p�P���(�u���:*"%��G ��I� �5� �8�3F���$�Y^U�ֲ�x?� ��2��N���!��-t|���A��Rx��h`�ucCƌxu�2�;�����]*8���C�뾪�:�����1�F��xZ�]��d�0wz�c�a�:��x툫k�/4?F�'\|���4�y���gN3�(!�(g�b��4��,ȼ0�#��f�vB6�q6#P����F�L�mį�G|#>�$��-M^׺�r8h�&�5LUPP�S���l&6�ʎ|go\���*+����<��ʝ��N'��8$�̍�N}՞�DP�OY3{]���S��,���8�w�-��46�9��+x<	c�k5˜RJO	Ďy	 jeU"�>U���,!<���1:�[H9��k��ZW7A��f�(Q�{�~������+��aH���o~��aMA������80����X��U��L��0��ȫ�Wb!x��[;l����#�!s��L��+� ���t�4�)M{�J�m�,�ЖBU�L�Bٝ4+}V<�{k�����5wKR��TߺY��D��<[����\�rx~�%��z��e�L%8�3�tS�Z�J|���Nˊ����_���;I�FJެ�b�t���UDF����4p+︫��%��]�W������%,L
ܣV���~-�ڔ��Kuk�^H.�v��aMy��x>�sNN\>���_g�Nc���M�8�ʒ�۩{�'�H`u�����v�/�ܷMʁO�&�t�d`-�$�/�Mt_pOv�N�'@7Jsgv�66�^�WlE-�0Eh�}P;M5�)CY�mm� ��-��;��kg�)Sp6��iW@�x�::�w���� ~^g[��߁�`�Z�z���Կ*��1��^\�D+O�ֱ�5�S<qP}ڽWu��j��������H@� �����K�u���ͅ�UD���h�w�7�&Y�"A�C�κ�6�6#~�$�� lg�x�.P��1!%<I��������Ę�څ��Z�M�\�j,��;��$��,�m�-� ��f�`�~_���������ͻ,��Dr�"��c�S<����!��Ef�n�������pB��ݪI�c���O
x���HRGx�'����$�������w��*��y>��ݭ�pjz���jy2�r��K��F{�|���o|���ۂ<?��������C�-#hɒ��h��A~XF���+��O�3��taN�=4yF9�<vG6��)�芨�_���&�V�X��O�Q]\چD��.dAH�[���=��[�;��U���a2սW.g��0�r��Y�Zz�G�ԑU%�;%Q�Ϧ�1~&6*��Y�̦��z
j$���r��_�<��i ���iY��FX|�������X(�����`Hz�Iox�yd��Q�i�We�F1�L���:��/s�FO�|3����}��cq���Z$�re��S?�m�[f�%�F%(η��]��<�����6r�3GRpmC�Hb}�-tN���d�n�,NZ��s��G��`���K��� 2�����+7�n=^U�Uc`�f�2/p�2�Mv�����#�k`��M'ZO�+�T���o�a�3����D��h6���*�V���߃��F��"DC�Pn
z[]��K�+��dgðĝy�������̉l�=SP]��0q��:Ɩ���ux�� ��l�6�m��z41]��9�=]�c��e��v>�&������O$S�VB�lXB�g"����U\=I�)�����F����v?yH���4z6a����x��/l6�Y����:~C�n�w���'�� [WEoދX�t�%�����F�4ӑ�|�����y.ʈ{FTc��P�Đ"�����թ^Jw*qވ�.�&�o�o�C�;��}��8�h�����$(��Շ�y4�MUr�jWK���Qh\w4��X�A��ұ]#fO�FJ6ɀ�m��8�[�ug��P)�=��U��M���_G{�Yɨ�Jl���W�#޶�������h|c��w�Ò�
�iwoU��~o�_ oh�'U�.==��M�>G+n8�+���y�������1P�̟1)�������k�����n�6}�$��a0q� $�4t�k�ïL4RP"���� l�'mZQ����BvP�l'3�d�M�]��<�Գ��w���ۜ$͍Ē��f<���#K	�r�D�a����K��{���)���Q�KE���r_1��$�����N@C�[1t�m/p�0 ��X�.x��!�c'�Uϒ�j �v ����V269Ê��wؗZo�r@���0;��Z��GH��Q����aĚ#�/�.��L?��.�+ ��A��@Nca$����sUh�������=I<�"��P_I��)L�i�t�ፍ]�;�$e<}��X&����g����-�P��k�T$�ۉ�CKeII��)xf}}��yn�J2��p?�%ݟ��ah>�P)H� �lw֊�Z��f}Iƅ5o�t���+��.�oiQ���Jl��!uF(�f�(g4�ߛq��F�	���M� �]Û�n�x��f���Y��OC�LGIj�
鵥���`����Rbw���S*0�r7���w��D�����j��e�W�,5�N̛sSm��-�vs��Bx_z��"��񻡗��?��Gc�b����vAbe�Лa:\6�B�+A�rJ?Y��g��I%DBs=�R�����_:cW���Vu�phP�uUd��'�jҖ�sx��[�F���_��_�1��-������v�`���W�i�y�/��.f�8��L�WIf-F��\	���}�����ճ��B�b��w�������)U�
ꝴ��:������d����v�_U�b_vBq.�$��M����?���R��ф]�>������(�]�+���/?8������2=PqE�����~Ve��g��+|���hvЦ�v��{�j̭���o��wa����G̘oS�
� ��9������xv�^�-�v�P��;�p4���Zؾ�ts�������:hnX`��$�w���v	eO�bC��0�GD��g]�*�r@�J���G��U)�P(� @�
N�뼞<F�����GN武֛\�z���5��u�_Z#�n;�L}�� �G��ӂ��I�=h_Zq[@�z6RF���|��etu��K�P���7"���WsF �l�jVc��n�YQ�X�[�6��(�7����9����Q7�^�,e��.�Qڕ���51��4 \�*�ӭ�������S&E����Ew�n�9/��Q��9�T ���N��+հr�򷑏��e;ӂ��8k&���2��e��U����o�=`�t�#`�A(s/m����	�BϡH*�5��+�H�(+L��o4{$P�z��c��6G���_}
R�����"Д?.g?���}�gĩ�����O��>�t}"p�R�w{g�V`^���:8l��۝�I�P�[�ʹ�J�i����"@���`�J���f,�L~��;����}���O�^�ז	^�q����o�W:�g�p��(�S��r!n��w�|��g�	��F���tuw��)���6�,��k}���8a�� ���2�5�c�`�k���L�T�`��Li'ƴv�����[u8̜�G�_k����A�#�Q��|�Q7B�nC5�H��K��_f�K^�?D�qG��{ή��R�ȑ�	���2�<��KwH:���mKJuM$�˦��~Au,�B)�t�a���~+:j�	.�o�8#\ďQ��j+��d�A��HdK�kC�9���(r��C��@�`��+�ј+;`�B�,�q\�H�R"�y�������Ғ��:T��R��i��R���]|�'R�V��ǽ����奊nZ�q�ڡ[A�Q{��*��pU*$��T3�.85�֫��y�d�kzȉ��8�vr9�W�m��n��K�l���k��رc�
�}���/~�֝ H+X�����ӭ���_�:[��e�[��ل���䔫y��P���kvn��hr��wqr���)\E)��}�}�w�s�kԫVL��cB@���cyߘ�?=Qy1k�GK���?s�r�"��<����s��MT~m��J�1hA�)R�Rm��O&��[�) ���>\��3f�h�A���8��ѐ�.-Z_wG�m�b?��5�Z���GDW`9��ф=r��[E:�@��VQ�ٴ`��i�v!O��X��R�Y�,Ʈ�Hr�F��������]��n�W�/�I ��vyqτ���8ЭP��`����0V� �F�1,*`���Y���m}M���n��!$NVL��+���P�0�Y�:�g��2�9��5*���%}^������אk!Hh��3��
�{�^�0C|�:��SD�j��8�N��M��t�����3��+w��.�������,���BV>�0p��v�>�v�����@v����0N��?z�sȡ�Gu���oH�0�#�)<D~�}�$����NW�Y�5�u�b)�	b- ���࠵�E&�'�}��iO���n/GcI�΋��2��9�șC���|O���Mjcי����D����iLlEܗC_���rpc�F����7}L��؋��Rț3Z��zfS�t�J����{)��&�x�{
�f|ÃÁd�Ć���w�	� ��PF������W�^���/��A���2@$�O��H���G�Ij�~ӻ~&NR���*��{1�0Lo.y����?E��hd��YI��{���/��A�o<��@V�V�W�hx�uZ�K�s�=7OO�؝.|�苾#k�
�Eѷ*ց[�´��O~��+��z
�ƢQ���f��A#��~k�M�L�N�mx�m���}m}����O�s*���]�����~?����l��H��Z�=�h�ݮ���F�2����\���Fj?��<����ڽ�j�@�>���s�S��lA�c؉��]��h=��d���qOS[ԽQN���1��P�Ͳ�:Jg����Y�0Wh��d�e�]WSU�U��B��%-��y�kT�fTu�Q�{5�5�Cb�;m`�d�t�e�]�B���Va��Fc�����!i��-S�Jq�?��X��|M3k�/�M�l�� 
R��aB	\�@��	`=6�0�����xq>[0�й�Е
P��3?�C,Ӵ`���H+K����v��΋%'��A�~�������r\X�c��BM�O�.I�j�C|g�mU"�C�M��-Ӈ��>�.�=�z䦐?��UiQm�
�!:׹�3�#��h��?��:�&�߼�ye�4i5�Q�D�I`7*�N7g����=!�:�$���� ��I�s .?v�
��[t�KwgOsE7����{i�U��!��+�NQ���.I��Ոw&�|4AS鏘_�d��&�Uֿ��_���;
D�,J����E�!���;�8���U|���;���J$u ���	{35)
<!�u����)h��\>���6pv���⍤�U�SK����P$w1��:B��rEXɚK�'/��y�ɂ8��i��(2\t�?��6�Ԛt�^�qiN_�݅�����%��w���74��S_�~��h�p��YAKŗ�m	�#N�B|Wv��˴8VEp���[׍Q�������L�"b�/ )�Q�4������az�oq�
�s0���Cf1� ��c4Pzw ���u����X��U#� -C�kOZ槤����OK�̵IͿ��ú��R���S#��&��.;us`|R�saT�z�4�'Ҋ�t�뽝#���vc�.��c���;Ջ����|�O/��h��NBP7*�L
���=`	?K,�#�R{:�W�2���x5�����I�t�Y����Վ5�6���7��\|��@,�:��Z�x��& =?[⟱�yb���5���w�*�"�t��: ��E�Ț�16l#\����?=չ�%�qc��B�J���%%����Bԕ�h�P�r7R���͹�o"P*v�S����{�XtN}�(Hi����"����gw���Z��y��P6G儹�9 �#�?���Y�}yt����!�