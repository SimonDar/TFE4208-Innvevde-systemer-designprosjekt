��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L��`������
�F���5'es�קZ���m̐�>\4T��Q����h�:H���GJ�?����@ni�n�O�N��ꮝz��F���;���h�s����j�i����6��J5m�]��.�N �g�XR�>�kG�(iv�p��3lf� !ǻ�7�ED����(���pK�Y��N��i�)ӹ��\��n%��.�}S�T�N��K<O*7RQ�@�u����D�u���x��$`��ʷ�$��%ܰ���FĂ���Y~/�z�.s��ON��I�Nuj�[$d�[kp(�>�YsM�"{���YV��O������#�˻ͨ�<ax;��.ҳ��io���\
���
�,�5�O~�n��kbti��5
�qwA��G��Tt�k(x���Լi�T:��+�1?N�e��=�`l2蹛�~4{`tB�sVſ���v��������O)�Z�������۲_�a��52+9���sD�1�fulN|��}�����W���~��g ��Ecΰ.�c�\	���q������~1Lj�Unf�:�?�#�1R2I�<�*���:�)hp��Q�:Vf��	r�E
]��+ќѻ�z�HA� O(n[1K�Ջ	�?�ߕv-��,�:kټ^�
D�NԬB)Q|��Zlo�������:,��W:�?2���8��00�����@���v�+�
����J�{�7�O�W�m,|L��:%���t���������ȝ�B�^w�@oӳc�֜.����Γ��2�'�JS ������RH7������{x��%E�q�#h�덝[�Ӭ��ӯ���.P�����*�����IR�|��%�#i�vYp�;�ޠ��=UR0X�D��.ic��QB�(-ʻ�2�U�K��㡸���� W��-�Ļ'�F�"X)z8>j�IO'��9�sY̳���BT�O�BlT�+TK�hK��<�4���.o���4�1�Ҷ!t�%ة�W hFv\Q(��n={N\H��^k̀/�U<�ɪ6T,BQ�ѿ���o��\�����#h�ߪ�wAF�@��~��U��-+�MO!�w�&������E�4���띫������$$<兕[��~_�
G�Y2/���/j�UP�A�5~�.Fs���W����� ��@+����&�.��^cv}��{�$Cv�h�$���	A�#��:B0�4�Z�aQ������kgz \�n�\{z`$��v�Y?p��`C1dwӋ��E".�h�;��\Na.������,>J�S�:�鈭����1X�r$sɳ}+�3S{�lꪓM��!��V�%��̟�i��z��gd�05�{]R[�j`����c��5ݜe8O�5�tE���=M,�/�s}?��RHC�Y%�A�H�ɒ-��1����l,G��{lvV%"&�|��y�\O��ڟ{w����ӃF�P�B]�RoX`�ձ��L=���s~���������k�rr:�JDml:2������_Tn����Rix���n����u	_"����u�ݘ8���6#
�U�����u�m�Uo3嫟9�+�����?nb�r�g�d�{���q1hk�:~.7��$�]V�Aͬ7�I�1���w�FU֜̀�E#� ���N����3��iDܨ�'������"��<��	��?�s��� ����,LYm��,��[��߷���
����i����C]�����?/���s�2ߢ�Z��I���<�u�����1�Â���Be�-�X}�˚f�*d-"Ba���3�$xQ~SS����v~(8��{'fG󯒦��@x;׀?u����\{;!�-��������Cg�0�X/�:]��e�o�z���eW6�(Zy�ǋ7t��=��I�d[�Tc.$�����/���^U͜�Sť�ƟՄE�}����~dG/�߶�'�q�#�l���Mٕ��3A�@zj���6,(���w�$7 i�/����dM�hօR�!�����>
���\� ��G\VDT���������]4e���m^�[.0�VX�7��i�T�$�cN��/�I���i W꡻}��j�+U�PZC6�����$��)��P�ؗ������Fz�^Ͻ봖[Ӭ�L��9�}t��e��=�k��e�;�35���Ps�2�:���̌q^!l���L�\=��-��(N���`���D��#<���U;G�#i����8�����DA����5���*K