-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BN+AZ5MSnEqhEm/9vFDDPnT0ZDKMXLH1NsoNMb51/o6ZkqberPp6huegWXaULjBXLKefBXQvC2C6
L2ym3sKzC951ht2RVyLTE50nMWzoUoKOmgVCruuo2PZPc1pVmiCzGmaDLdc5MO6dgJNAHVDTIxA/
/WeN+UNGX+TRt1Civg6/II8tkQMIHl3FvwSTB6gPkPCStqHxYWiN73fck0sutyObGrgH+gkwWWlG
Q8m4gcAEEL/D8VRCArKAjE3/LtRRe72Hmmey3O438XfG8qz41rQEuVuuG/ORrJ9zVWD15X6zKxwe
s6ugy75NRd6LSPYUIrjCPPUzKCLyvtqqL24T+A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
fHG5XRXGbgqd6v6cU1MaZf/D5ajgbIRyKlD/OB+zExGnv2STYwBShz6XmUoaBEe829NAxnbof92D
dKiohC96fAMH1F0t2ZAYWQ0pCshTVrvJnKyLrd7OzNjQ/V6/Qce1byn+OeFmss9IWVt/ZB8m60T3
RkNk2FMtMRZhAIkkd7b2utwXAcndcec8v6e0OXuaeUs/kbmDxb6kunPEuN6npJmPmv1Qrit08d1Y
hUAZ4ciCiXbS0ACwilwUEk2phnYjatnpdxLQ0r01wQR+JmmAvXok0FX8tg8hd9tbo4Tli88/n9OB
C/6NInU695JCrj2WdpikGq2mhY0AOEI/vH/AJ0I5Ahw8Ju5OxLNDvQPnKXKUe6ZYjp75pMLbbqNk
iVqRO/Vz5JpAddq+NaGM9cmyCJKrSa5tYPTEdWERH5OlOWZMgDhdIkzFJoIsPxn2xHQwq9mLIoxV
2ebRDX6/4N3pEcxsq8I3utlKKfM0PMIDq2gDqZESsyZUzDb0QMA0lAwh3Lq0waWKd+iPNS9jalh8
NorsNY0qlT6ePXK3pC66WH5vifkb4/rjrneP2R1D+OmZYCa9YsYjEePcz0WVY/xSD/DPNbaqEpPm
9Ke/4z0Gm4MecqUSmt9FGi7m15CFrxUBvFd3EL0cjdR3e3aP4AiY4gGh/1aaA71z+rLpDWdaHmVo
5mYqvc0Zww71/LAhSzP+nNJf9SQYtA8IwOt6xg46vde9SIgJKSYEaniWmfcsE9QiHYF7/z+jdx55
OXQqY2TMbNYwM9mkCiYc8mHUREGnQPOyfRehQLx6gSPo6ZGKDkNOUEUXHCle7Xmt9/5veqEgKZ39
wqL00jCiK1ssmwAWyFDrK9AhXdZxzS+R6XA2Zsb0X+WWs59GWucPXhMZ2AfTdIN/NETMYgTjcBAu
Ru8evgYs1SsRDKUD+e5Gl9IW7jqbPPWyx1/X9ScAzfYrk5MzgBk0v1WQCU2xPzUXpmK/TqFvFZB5
+sVReEO+MY48xqjjS0k9U7bLr0GkqDXnTWnh3diOGDZuAg6QHCWZbwdLUU9jPOrFTNs6clDo9q6k
N+927Lq3ULOk62ZWn0mB68tGVtk9ihDkjBXnmDCThfeeUIh7pPwOlfmbwxnZelE44T7Zlv00aN7w
XwJ4qi9cXs3lOlU4E50x2ViiOGWbAAOEhQ3DDSYxs4HBgFZTVdGtQ5r99tCYv0Xr8UZBlHmaZiOh
ak6vp9+al8yTeOZeN3d1z4NRmbvkVv1kMVPyzbPtcv8sYmDYhguuukNCWT04yXUbnENlsgorzmdB
8ugREJodnnycZ5slUWf6FFX1c5zjUZBXF09UyYyjlLyTUkutXQZdpOs9QZPGdlBpem2M7jvPZpTv
2lEYgQ/RHind5qbIRaGJNcAgGmOlOzGivTuIKZLKO56mU9fORUKgDwCWiFxpaSo+lLodWkO+ASwb
imTsXEugNFJliaKefNMm4mL6GC12CJxIrqLEONl2Jr/GPP2o0ex+gebzkQtJPaPRYf3pbeluVlVc
/0JXlUjh7mE+Qx5rpbxNiiw5DGjEb4jX+SY73rtrLl5Fsl2xdPIJ20yw19BbYyUFU36dmUJWP8L3
/7R4rd9W1ObwH1bh9G/j12Pryul0yHd2WR2uI4LTPgFTZevKjnCYyswehPOpqdUtf1mG4koH7zqt
RL2Cq9G5OUtFkD/U22rZkk4tnAtPBpjlhxyymGfgmjKpSzUEeeKXAZLxgg3r/rNHvZHx0QGI+S0a
LBQbWw9uB1rO5h1TsdvUOQ2xtU27lAk10ZzBR6tkLZ2pLHfuQv983ltNorc4Tw4Qf7LvLwObPinx
jayMtQrYO7/ljOaTbPDtwwzOyNruVFFROUKotKxRo+s7ZcKQ6JzViBiALzvcZjF7iYLSG03rFMLG
z5hbmWGUiLJHT3gDiGmWC6cxfvHSbLvglGppYByEdaGh0F8KruLR2rKtmlnSNuncRfPl+8JjBC0h
qp8PGseVc7eGF3UWx6uMFCMFWqSyknEnCdFV+4sFIU4TxpFXhJ2t++BhFxvgF5i7SEamAW1R0v8z
S8Yg9YeWOg7g5oy534C1xvlu5i6QXTQoDn3hrqRJPi4Ee3aiIoDaMRuQtERR+R2vbqMd6hDWxqXw
ZSC/91zvxQn4Q8WNg//iw8SJzb3bSRfskDW6RpuGPzLrA34qnkTLrmQ0rA6Cp7Lp/lRspbJoA42Y
c30CZuzaBCI3Xb9PQ+JJLD3ij7lWj7C9GE5mldq1a/5XP5TMbGDH1kIDfKEosRU4YHSDVhswcEnG
biTrn79aE0wBQfOHC63O4b/owEj//O+4ec1+23E/7s613rSkUcVSjiPDeKtjy1xP5rOtqlTVSbhb
8gFHQQeSJ1aHzaykZvtUMebIgZEZQeXdzYpdx3kQkMzkjYTO0cHXka1eAeo5oxNcQpi64uNARW/7
MAq2HXj7S7jawvxnODELBWWckbmwZf7g2G8zZQ23XYKQDCvsVoSjUfzV28smMjsmaiKHgK28glVD
RBdAnkvLGniE/OsG1mrwGGAUdF6PviPP7zZ6WGUp5HaUTZSo8ahcdqk6IB4S8zZAarsg0qVtMJSq
/qHyVpc7QMIlNOMmZ1r80AEE3C956QGky+uYYs2GutaGtdHOJ8ZjyhMzoI9PAOslERm8Jn9iCceJ
2AyJ9E/nxP4xCL5xYsPjVSsVfwvOfcV8hT5OuHqoUrFXYhQ1oeCrvrj+gP9o6xxRZG0QYMILduUI
hCItOKvzPff7NRXh7oTVShZYtW4GHTi8O0jenkEdbJgMypjQho2RAKzwutw5SbBw+ijR6mhd1N8H
atnDG/HxMydAT4NLrxr6vWvA9MlPFBgIZKWCyWmSZuWdvF8B13At+mJyQc7E+2iw4E9Otql2G0V6
LT/gsmB7/5SKSe6yoPrpJBSHZJ5VvtofTyDDKCXbzrXui6KFz3U96Ah7kOiYqG/mt18OKPHtKtcd
vGOF/bYjSFf0j20Nsao38L8JD+V1C5SU+neqaLqiI9fBUTCGmUpNrYXOj/qVtE8kdvCvY7whPMWw
0VV1O02iPbp6GEG08plCxBT0aeMfxNPm/0xmPADyVw9NDGeBhuzJbdi11KH+nwEZ/ktGUbA8HRtu
f9xK13SniTL6/i0rAsuMIfXJ8qkxI9JM3zsdWMmVUJXrKudSXSo1Ba7wZJBr2G9qFMUdxhN4VJJw
ZzLDFgdhzKJfbKvXZb8rxFHG7SOfYw51oqdnhwX0kZ24O1XssKrnI8M/jYXc2lAftXKycsA7ia+l
t8WoW6yIrNv4gDbgs4i2au7HJiHajdZf0yO74kz42REbw8paVn+VTRghfRq6ObfIeu7oxHmqvX5L
ITEgav2e+ZC6jsHRBuNP/gzPuI/BM/bNmya7U9wOjCd8OBB1aKfNG0RkUs8m7Hg+vlU9JcqhUVXp
RKwfx6B+7p8iJ6sLQaSk4gYdfsNmNHHuaUNYTCtxUfGBEsdX3zOgwXCT7tpIGlMpT8ubKN5T8TQd
JXyK35iPK1lqvK+szs7eO5tfvkuUIADwLnoJhLu2TfjiYzAn+OEeclmQj1fZ3rFPIKqa7qn9cktX
TERSYerPw0aCzMaYQ/Jp8n9Solx/CwPOfEj5uppCqb52+gE4n+hVuuzT9f4YWqWedyT88WXOez5U
KVv6l9ZmqAjc+u52cqGvzJadvDh1VMmMV+hvjUITblWh1buWvf2uddIj8D4I+Wrp0dncxncXq61T
PO5/YIpGodNPegAOmfq3xh1YiDLVIV7FtjbdYzokP0PjzGxwAl5JQx9b13GtBPSlxB4pC0fct1cg
cj8FWKXI9Rx2v9tOY9kX8rrLbkVEp3Zmvw7mQj3UrxNQF8uupDfyiFrNELW4rivaeRSOfqXaW8oj
nyZWgIyFpbNoAnBgq5Y+HCLT9JPtBslSfsKveLuAWof+XjMKtv/o7yCCJN8ypi6ko2sYL4uvbI1E
B5kkUBevHNT3BXUL3Xd59q0RFDJBFnlpDSKJ+Esx4Hsg1DBMWiXkjW515lxmnGh73Z3TgK48wnij
DHd+vSE4wwJyFlGiC1sstMpCFvp4IlrE8+N7XWjzyTxMr6o0PxI4BC60LKCzPWPP0PaRTcqOXYvh
GKSudFalGq42em0lhwhVzRo00jn/9/dGMOO1N4TFoRbax1XJ45HYaXjgXB1BFbZCRksnKSD2xmXj
AO1LhNMbb/NkPZv7HJQZ+HmgAxWZFOKeijgHODyivEhJrDxLMWD1URprAqQSzTijo6G7lO8QSizS
zjV6g/fPd7yjHEezDOai77MCFvsGqxmuOYKOysydG7aPBScJbOQSNakjjIHtsRuAlhE1/oDWHlNl
olnBGUXnxgnKZLUY6sjeQYLv5nEOHQ4N86727+cv992NVB/HCzwGzWj3z0N6kRRFshDUdveOBhGb
9ttTIDMAMBlNgM4Fhrs2VbQTDDnYy4HK++kRHtAxFNwFh2Hm6EmgGZGZs5VwoKOaGZ4Vxk5/kwMx
8k3O2enlW6G3vAh+7LGyezY8pXzD8B7FBo0JgT6iixsGgTEHQzm0nLgHqfPUUIHzNn40utNti1So
pUqnE3YYHRVaTvQ/liknJ7IkDQM8ed10rwAfi7AjFwrI752z4X0tlifSaYPuinayiATKfolUImbm
Yw/nitVakm1TMADm4hkA5wY3kphtJHmxvfhMl6w0o5GzavQDsmxToR+SbOG1yNrbesQWrH/NvT+U
fY2ycTdwyZls1RAneFSU8j33abUda5LwTgdgqriGu1Peefi+QMlD8dcN7RjC6fru5jIjy7iFTzbN
C5sFeI6HmKoDpDjITCHszUhgyhs68v2UhPE7Piwu2mmbQsr7ZINHuAg+8cyaOGInlfZeYWlGAmcV
auXWNVV+3LPg7kY9e3Xz9+LSAhp86aIztT7zE/WbLPuVvZp5fZ/l1LiSZfV9XB6eL3mIatSa6XFj
uIlRUAnmEJ9ZfDTgEw4HLpxEwDiTAjBct/+GQm9wv5itfrB3yWWCJeU6iXlcUPGSKpHyKbZYnpUr
7kCUAkztrkTsCH0QYUhDgsWxdFNXecX4JSsMD0uWigTqIsuYPo4xM+suvNJsQhunkV3gGrdBT92i
3AHmmWWPpvnWcY63TL2XPBchMCyYICLd/3lByQG+onUFNNUDLKMZ83QqFe0A0ESlMLT0K1O5aLB2
k3+saRSzwGaPVRqULWBRzsxKTJ8dpJVul0nxAJcE0XLofmYziphYPlje44IncXcmn7XZkRuoWDxG
1tyTkXIenQjXcaSUYlCSZx6TqrG+Vv4jcZD/sI+Z2u66ij0P/9i5d7Ns0KmogXqQJra0oOJ44GoZ
+fwJmVzG6mj2tzOZd7xTU0DZ1CZZNjZvMNe+QNZbyrYpfVyOP6RAOXsT/BJX62h1L5YL4yL9Ezk4
1PU2p+dPH2ZmtK/xRtZVIJ9gHqb4p/lWxyFAyu8eP4tZ+CBY5iC6LRKzzKp9AukZYNYLQpbvw+iH
k5VMLRX+XrEd6W6rHoscYhz8KQIX7jKYUG+41WVcA4IJ8RDG9jlEvxfjKbZD3xjGMdx2FKIx5pxg
mw00IT1rcwA1064mHmBku6X2wiEJ0L2KNd7gUfWWYHdPS9KYxYxTJUTpZOE8vBTBiyikm1s2i/Ox
LllrAfcQL9v2ghdiIN1OXmrE739tRc1p2O9L8v8quKw5YKv3zfSrbsCoUrxyrQOLD9FH497zjoPv
PRLEu3GrfxBgYj+30FKu7bZRXzO1Rn5qdEhzaIYTqdatUUD95JXPCrgEIHMyIak2kgWWA68jiWjz
Dt2t4aIDBEJvC4+/AFlNdaz7KwNOzJtkqsBP9UZuPKMrjjuDlpZnttZrpW4M36tsCXxFR6MeJIbS
VsJTshdKWhH2V2X+jRtKtL1n+uTplfQt54VcZawhsxq8G9X2mmrkE/9O8mBoEqp/8cDIHxvXZw8L
db1CKy5RwWvrr8I30OTB0UsVbS9Hptcnfb4SLRHNoR2II0hEDDT8FJAgBcy3XoaaGCco4k6XXH58
BnwUPdC9vtNCAaMhqu7teYBKTzXbuBf+15Mg9Cl7xvpUi8WnoXVSSK2OHjZ6bU27kT4WTe5QMiDT
3PWkCkaSFyX6xo3c5Q7dD+w/sqSELBU8mS1M7lnAEjt4IBS4cJfJHE8C9BDyrBq+wjVcN+HJw6qm
UI66jtJeg8IghcxwoiKU14L6qrg4f/vqoTjv0f/fwqpUPxZXUFzxqkLiXwpxVc3AEgPhCHeoyk57
B08T3UwfANCKO9oHq05p38mBD+pUdZzeGd26gb2rZrWvM4nn6TiiLxR/5RyDuC6JmKXpSvVWas/+
bHtyFCfyTsrS9LNlPYk/I1uiKCltk8HHYWlhX8p588X+17Db4HoOY1qC5jSR8qdprBZtrVTCw0Oe
WXnfb+qXyvkOg0Wq6J2WeJk4hHilq6nRbqWcNeI5JPbHj/f24pzrncMO2nl4zT97x8WWPaOCIkYA
09KZXPK74qrgMP532EkTdx5/IuyZOuitoFzL8RcmzO6rOO6pnxXshJrKxOh8xR279emoDumi4sWM
2Z+pRB2YE22DF5Fyr79125EErNx3e0mq9C5P65wOBFHUK8fg0oGBjo4H6SlChfZKeAiJoJ2G6IHI
I10Q3AUpxy9vYZnGikehOTNjKEBomdhUk3MQvMj45LAIUzRlrGBC5/DQkGClycc8a9CmfKKz5m3D
8SUdidIj8u43Nc4aZVCwzw/YJjpMCaDtZFbIrP/XekzRRA1xAdRDBNBoc7giTQPnVjSLMgLzQV/I
lYJnnxz/PIVeq9LeUFj95VahXHlZ/WwhvIuc4V7t3MwuBo+WaedPypKuMeJRCrSw7kRTz9tV/cww
lFE01sXZbifcgM2poGPmwyGNp6yt+HNHLJ4an1dLEaqRslFUgf6wbLeBpaJ3rhjIsJ963QMOnS3Q
LBaWQbiXCNYHX/cBum/4qpsDmzI+4Er0gB6yg6tidFD44TAEz3+GOoSLnRQs1RovjdogLpZuXxqE
wirqNWGjpiMnEyQwT65d8xLKiSOtnY/H/DWiy3k9+izDuin6jTPYRSRAJpdwGezKzleAOd08/FDL
I8JXHfKzOcqc0HagIg8VjZUJ5mL4G33cmMTmfJDBBeP7E3eMVbNfaSrkKhVyGVEmG6s9GJWdmBr6
wxeTEM07Jh5a7Zv6pupR/5x/NL/bTt9NgclHVjLfAhlDJQ+/yqBabO8Ezohi8n26eSV+FYH0LS0c
ak3xFZ9Y7FU//KTEaAqwsYY0uVinvUckso+KKNAZobWQIiiu1dLUPOssgCs+VKF2udQQ/PFJds5l
W5RwzMoVdUSCfoWtISUz4qUfELKNtQwYpo0QMvYqMNwx1pHvvnRuPDUvtGrO1WhdIcXq7KYRphXI
4w1DQOGfA8QSex8sQvLjhdys2LBrTT79uxBlEbhjLPw96yhKdpvwZSSrznDuyr/u/mUSjf5xucs+
f4+HF2N6lsrp3VMrKzcPWsdrs2wbs+j4DGgRFYSFVQWkjII5y64N9Wn54DHyF6bzccZduvntJ7x7
ehgQjOhF98Y5zToKLUcCpJbIi10VOdglh9RsIckDd7EzyhKNgpAS1A/FyXqbFxcpVDLnUmhnRbXQ
1eIzymsjrK32+n5Bzhp/2yqHPyOdD6PHKbP3Ut27pCTGLXWzOSJW1Bh8qyQfyjUSaDikG7vxWBoe
YRBrG1iO5dsnunkjUarqPyNN1gOZFSNGMX8FYDId7hfr5OhYJ9ssD7DAfQZKTiit3KCmIDF4ktWc
k40Y9RupEn7b1dODyCYLOA9JPPaHBy5qk09EpuIXWjQLULLBAz1Vl9//5LhvfwHMFAoboOmsQNLT
kdqmCUDWmQHv8c31WCY66a0kK/CMu+EtuBk74tnw6IXx6eiwADMyMMaweAiH2fHhZZXpH8VuxxJl
CAeZYjk+0nqU6Hi8ixLMXpzwOsiiQsfuf1ms70xqpxdd8SGUo4aFYA592cbZlQodXMrdeVl3WCUm
gPYi/t9Pav4YIo9giZonE2CvIIyPtR53jDGTwPU9NTF7Q0w03RP8jgd8fPKJSye1dqt88leZMsWh
flKPo8Gvsbt2Q4tTvakIAVowVuTmZTOI5uvG/QRGoB/UzDwHCyN4g3J1E9amlIbkJ9DY8d43S2qU
ibn9otgfT4QZGcJPC/cDOXYIXEvTVNTCV1b7E/zRJUqILgLKduBRomwBPm7HGl8vR2i+a4RpNHr8
gzJo5qZDoYih3gQ1GLSlsd/UH7ynNwI82jVBzSxqkHX5um/shY3h85aPpLgev6efVLkADdEyeNox
7VJgEQPxkXKU+VEPDszAczmhLfgBmwVaTEwpO+OHAyNRlWs6uXc2KZXDuWx3gMhGh+ppsPCBLK+f
kG4CzyKdYrwOk836q8BTMt5/syvot4322gx297DrnEhskrq8kspWLY+T00YAhg1txqWU25QQuI9h
9vh0EjR96i4ftJ1im6ZqasSgUYqiKeMWzpWBVeDyhbgUh9M1z+49J2ql4vSL5c1rlA35lhmXXePg
GSMBP+IRWWJ2TqAwD50rZbrWvpzWJ8C/yQ4MJs+hObDG184msRo3AoVYEQAf6E7n79fFO58e8TVJ
lqn5iB6V99k3+eazytqsWEG6XaJ/7sSurmNrc88kgrnvOVOzXKHmpob6FGdLwyyUIjTJc9T1FxIr
9SvMrWX7GfDLYgHw8EyOf7Knf91P5RGBWgwYbI0XCIKaxuDE1BjQJqaWBxA8cG+AuiObsqqPwqsn
4DMBlvgb4KLWnAmXxzwbXOmtJ2tZ3vh10etbUESRjhdYVDB8R25qda0t8EV9aLLB9hLM0v/j+aaM
QA62ouwWLDs65H3JD0/KTft7sg0lqAYKEDuCld1Alyylw5IqtMibd/lmcj3Klq21wjDcFOCexqsU
odn+CJDivawt02n4dzEkg/oaEgLJnpG4TXaK+XJXn8sTCGRfBxYw42QKne7bbIcXiFbthtD3E1tm
07U8fysBYuKRqtUU5COe+olnwUyuruuEtB1Il3wSfwh3E7EYovxuzwbjo/Vcm8CyY+iY6aSTd3Zu
61T6htbGLetquQiusYTz2J5wBghUSOA7aTrZC/OONqeaJxXcs7whKkem4zBt8sSmT5onLV9eOFW8
y7UhJJDFnf/IQBKXlzb9/cuIVvYYUadNkgyb3nS2Qt7/5SyxoXx/GmJpsrINSFG4HPmJvlVmV6z+
l1dY/XxYzQ0Gj7Q/bzF9auMjd8tSccOSFDa52s0k9KDddEUWQ/WxqCM4ycN/RPm/VaJnlTTbgtOf
wVH6Go8IC+lMisfP1r8Se8zfXd8VvoKJ7WS2iK/bs1r8C5+TnpoSaekOE6mRzSRMb4W+yhIw2+a/
/h5sWfX5qyxzPocAQhCKAHQw6gS/eptDo2quhoB4QVdvtUuzdwvwS5DRp3UbEF2uCXouOi+3oet/
pyL/Y+7TKOOrdrPusBye8T5V6C9F5hILO15mnORkXlicIUoj3VkGouXiSq3qgSpNOzN7ix4JdVCU
wCxQusW1P0AwNoN3sf07btWVM6E8i2xFNTOA7gasteCU/I24UzjrnqvI4ab7O94iSHSrak92j0u9
hho1VHb+xW7ladK59L45dx3YQgIzps5rKYyr3PRjrct2FuPQuS/OW6OYKonDgATMER1wPzY1ar1Q
hm/dMiAv99WJJWv9wUQG+BDlb/GzOnu/yShx7Xwxf+6gbnojh0fO/kl9I7sjwCpgACkj0Oc6Pk/o
w56zFFrsskRyIeNASZNqRgG1ZlTgc2adNCZqN/dcXifK57JVDqLi81y8DsUVwnyfWNosGtFYFBD7
Mm4rCscwD0w3tAznZWz/WUBHhzQ0qEDAO+fiGC39rA4IlEO6IwBPg/uxHDG1dBP31LI0uIclVwt+
TBC/S/9htWARLe1n3fmAHPyNaN33pfjerhW73gzfw8yWL1AVliQ6ImpiDYjjxaeJjcsqJFmn0Ibl
os4yD1ELg0kOr1QOoJ3eMtJnpfhsQBLxCEImRXjMbCQ6n+LDdDu/GGEPNGwoSKc52prfrtSF6SMJ
/0MFCsa7NJuZtT6xo9e4dnkvGgrxJucfww2A5AQ6EYoOo4FPTOwmd+eGRL3wePT3BpyFymZHw+sO
Ju72kHwWN9SkGezwfFAHxAYRh6zoq70kOrtnqs5UhZiwRGn+pu6xh78HbkUKJS5yoCebwTVPD/dz
L0voavEba/7ygKS/cBUe/yA62FReg1UWWAMD0yXcEyF8n7Vp0JQd0IC6E9nj8EfB4QjBiZUBw3o+
TvD36WQaKpK4SnhSCEdNqO3LNtnsNZ+VT66JJJrBRzJd4z+Rik5lv0j+DP9AX4cntDU9zKMyjsTI
Iu3G8x5AnX8eUTh1mQ+55uZJKXOQ+Tv/XELeXt/2EblvSE6MYDUK8RcHv7NeZLacEiMP1xfcwmrP
EMzfkQbapnwJ/M1++XkAO+qm4qtFQv11L0pSCmtjkYOvlUk5bcQ/BSsqjXibPR6xqg/NicJpj2qh
HAzNYm92JvSyg6gic9Fch6HGk0FZlV37lGhFa/McXhkrw+LZQtvxs27wX/HmeGjc8EDU2KOC4mRA
ny7KPDzsmJgsPeM8IUFGB2YhjDEDqWX+pkybksVL2Ca/eLJI0JJM+LDhc/y/WuIZs0DpzhdOgOut
mAt3DPu7DHbl8nTQhnSFGIm3SCUsNgMU7KdZnTiOXZf0t9VavaZsvhlcSZwssl7b2WwwdUm8AtX/
Qm12f0WyYmilhGD5n6dQyl7bmIorEZMmkLjp2xg717+MRctR30F0iYdVVIldusXtJ1Os5ys8OQ53
JI6wI9U/b0Ifel4k3LX8JdEzr4bsIoZ3nKg+z8+EpHtxUOHuxlDx7PJ3Mq0oLVIyw2BvpWNKe1l/
Ne3SxStzvkLo97MnEsU1nuofPqyfU1O8TGuw/k+yGpjpNp7av7lqaZLYvvm0desbP1/wfi4hYMhk
5D9vJNPRDyQI9RQbqlTd+JrocKWPia75D6K9heX2kSUsNyOGn+oJxB8r8WUhPxk3Wm9QPkOTQWQf
xo8oKjfpnQ2FkNNSys/P5eTRueIjtyg8tpJYgZP5II0djPHlRhLc5Pww7mjW0jZPTiKyp7mVn2El
O3o9eBciJssJ9Lh3i9Q3sgHLo2ggwKXIJMMZrO2ZB55vV0hOpvQ9KTTB8sjwt8vm2c8MVAJjn8go
3Zxnem0h/DbpOxMCgnVjISa4CWN9AuOkhf/ihalubLx1vq2GK7jz2na17iBVNgmj2EiJJ5uyTV/Z
lclQj/4iyIX+TBqLtxuKjphaPa6G87Ig4P9mKpvD5hfHWivbCX9eCWavpssCHRTbfv9KD4hFmTET
COClmuzeev9YCR4nKNRh1aQLtWY6a1D21SkfUNlrvKrShrRwIjvYcPp00YQFtmgVW14Hg6wfROT5
76zFFtlg/CteEs7jMvP/ErXMJF3gCDpLSU8E52EVvAOrGL0CHb+v5XuVHsjKQIDfi+tR1zuKrvHk
8YPmlu1mjv1iK3gJ5c9Pp4+ltMEZnwEJ1qD7IgeMA9HfWPbpzalVdbG/gZ5s4WteJZi3TePHB5sK
Uw4S4Gle5oVC2KE26AuFqKnukCkRGj1u6QZDWobZhopPnQrm79dHLSlxRwHPNxL8uqYf9l1qWC12
zBKKL/mdUig+Rm8y+c4QgORxqQExsA2FzD5uv1inn0AdFnHpEh7jSBwm3OLeAra3FbTh9W3M3VNu
sU9OdFkHacObYSTkd57p0Tr7XlvJ3zoP33kod3oicCOYIG/95kiGK0BB6NciZ1vUXYLjHp5b0X+u
GEPWR2M5BIbKGkCWB6J0bCGDYgNxFEm0AF+Ks9xM7YP4uXWoeAdMt8AscDXu7WJ6ttI07T7bGtym
kOjJKvMrfOn9FbzqkHHcPmRBRFX1vpmm+azH3WzoFYWOcf0UkW7NPmJzkj3uBtCPsJzuOwHNLpND
b5rkBQSJnoT4ZFCe/zYceQXW24C1aXWvYvigfGU8MNbYdieDmayFNribY/16QS4c6eM5/OJI+DPB
P72XnSAnBIGlW3YB+LJ7TgWBhX8Cvi5F6AyYRBDsxigMguwk5Uu63uLuCnV2PFWd8j8gdt3LuEQv
p3UOkpI2YiL5vqXBiMOTPrAm7KsNCHCzioQuNOj+nqcYwP1rY7ijtlGmHXY3hqoSr4QvBjknfdCX
vZOeEC+w6cN1c8kcvBgEcnfSbWdMbOXPUOvTZQmlV2jpRydftQrVaKVFKFHM515PGtuBY6ZAXYDb
xUMuLyLPShp1QQzoMiyZYZ1X+PeZRkYQHT4cYccqC02YB/VMbGV3Xmx2SrHWDOYwUym843DKiOCH
z08yU6UzTlKonTWBHD6AdazYUMqVdXK3ZLtjb061MZYgwMWN0b3Z+oXUIJDEOyYljlGHVWguzDCL
CPgeUedkYlnxNvLR0gLeH42tUM7doVtlCPJ/Qr260HrO0xuVBdyntyZysxlSFssGXwQ4Cjgxozd3
b8PDy78LgvDz6hVNcwJyR0BRFEWZp7bPA+904eMHSVQqEMu2LkhuqgNzxICQKtXLgFI3aiDVR8CI
68oJGwqXnq59+L9yjJdMi9XDpo1QdoL2YzHDAr2ASY8R3LwYURIsWxCBFprMsP2CZ6XhTpEspR/d
vNiZWjeG0+s2czoYpX4ULXZfxoRtV11ljkdnFTFzz+DsIOo12NivkIpvEcCLHzGtvQxwGtxQOTya
V8XPnqQkVY/GV+k3iUYX1VWof7GQzjKAJ0XbblAIJ4LNArpywINL2XA+q3UrSJyX2zCVf6oC21MG
Qib2wIlDisRnV5RIdIgbOM+m+MpRfgkzVFD9zk/XNgZ1VrDMLNEV0Me+I7TaYqnI9lYqlON/3RoJ
BggT4CkTyk3oJWnGNVG8JR4HsAqFKa94KeZbPe1/yQzJkAw/Es7RzLfG2sVw7e3x2WBGJkn60NbF
4zGUC9HLloDrj5y9WkNhOEycg5CrCve80zKu2oZb13BgdMC0QJknwLDN5orHXErnS4/GmxHKwfZD
kVK54oATQhW36thify+LmIhYpkBf6sljU1jmVyCq6Af0kVXg6P7bhT7aWKLsm+CCD32KCDRDqzrH
0mHOm6wBLvw3yN/JZ2Fuo5tuZXi2EVOPp22p8bZ+lt7qUdaFsh3AEpM1IClx7OFei7HmPtiC/nzT
Ji5YdTRbGTH9gyDMZv9wGyphSGcJqKxoenzmhwB5ufPwmrzEv48tuLga9s+cl9UoNkPZXlvzVZLz
fPno9DbIKso39e6fbHqFSHt9a58E9fqbZLJGdrPtJLziF9+GyU3eTVgLJWaZ7MFqqcWMK+j4vKxB
1uxKk9yUuO95OzR2WSr5lZvgsy1+abIZHHEOi7va8Az5sycsA3FazgFA2HvU1Yw0pn0KI00+s+kQ
OBWNsvyyG2J+oIoGI8OmgpCrMmwpDPFiH59pKFTUQQ5Gtf27g5rDVPSnXnf7dae+kIKjviA3MNFG
JHTsMLo/dYzs695Pp4+kp4F7gQpuqyW3ZTD45cf/oLHDJVZlsvZ+yQ9Ddfwqy59EQB/MSvtidcZo
+exW1tLA7L4ldEe/8LtmDOy3GV8RAK/k6FQ4uyMckhrnpwA/xtQrJjFCZHooQPeGIIrxBy6s+LXn
3aaUSqX7f6KA2jwDomXDESD92vcHrzkZa8stSx0mDKl2S1TtM1NIYQRuGbGlx2kPmnvvxmfBxfA/
wt1QDKFe0rgrXU42CJEyKM9H9D6vdQajlvXBSFlTE3Ba4HneFVXgH4TNgOooTwNgLDhUsGkVDGwf
OiJW7GuAY7OISFCQRz5t3jfCZ53/pT/lrFt2w/dTFietLC92aMtunOm7ArPSuYjwra1Icd8KcAt5
RkWX9E7sPvK3fSOYHW4bv4t5Y5PPvm9jo7HPk/8fSAM36Z04FH/2Y7QASqAVx+tD3lTw0vQkJzB0
L3Rb0NTGGkMBNcV0ajHVT0ogWp4L3ocjlk93VQtHJbMVoCWzyv1v2uCsvwdOj2Hiq2DUR0LTNUFA
dPZ/nwaPfmfrbckSUnsUqf5d8LMqdqpjYyuzx41l+zRm6UyytRgRLK/y6bfjx34fmvhyW9Xy5qmk
0WbPaHCtNau1gRPIzmit0iRT2NCh5Ha2UHq/Vbt51tLHnIu7pqcSZZEUsYH0I6FoOLSHiDm3yyAb
KlDUpU82X+//f4DDgwg4EfcFvzPIPC0MPOtJ28pVd1FEgTRa/A4yvfLWBv2X5qelndTthQBy3iCt
o+nUTmoPAX6kRudCypZWIobXy1G6BYff5Y5TQCimyY50viFFifwW5ZumiRvDgTP4boa5zGpVT+II
n1lef2NEA9xjWgGdaFiwq64mT7AUup8jlt9zOpAdGXcjIi/QWc5G25vITUsrmP8JAC7Ti1Mdcz2+
v7OryQO8AJbd1vLhLX5UpM9lvXLLS5ilXDxpeKBXSZ3O2TNnw90/t2Jrd+U9G/xa0FC3KgGngvnd
LSimdHoR+nskL6EUl7QZFoQfRw26D1FSIv7eRxYbvyxR6DAD+gsZtDcvCfSsn8PZ2gLGiAAVOGHK
8cs886yBBTJfiXMF9h+TWThU9Yt293uRA+n98A0s2tQyKz77HZl2QDt6fTErUFc6CVfxdv2QkHo4
4AN+mKLXK8iLI3QlNgtuM4MyfffRdtVAwixz/xTnjIokPOmcKi52H0PbQ8B5xeJkdvNOpp4NvoYQ
YxfyF4sY0aWEptHEgSyN+k5OWe8oMOfoRCpDG6OxAg97fdfBjd88t2cIczqQBgZTn0LTM43h4Tvq
5n1iXIEjO4c3ww+/A1iLedo1EN0l5A4eyo3MZ1I5TrpMMmJcbYPqfpzICXGGm0SjZJXPWvWo7Jtj
fn7ssZeWuomt5xuwxSOElp+5Y9GDIHNr4ZgMq1AjAw/tFUHllYSSUeORjivaSu+UDLZh/KQrnmOK
Yo6CZxp1KABjLCapjPQDU/9CZF0TUGVB+ndvEEnv/fhuNixLqRiX8dtKtxQbF8vNmlgmB0ZOWBe3
d1ohynA0v7N5UzTELS4WcSPn//NIwLyjY5dD545W8N1ASSMbfwxunkmxNC/KoU3UhKlX/02q4jrH
j3CdNG+UK2J2jgBUIgXR60ZxhTJ4WIelMomyfJU8YfVrsTlYX5ub3XBW0OAA9A8ijAsIS5KKx69u
R2nqMz7yP0g4ah8ViJZ1bCfzYyGi5xRNwWrlzj4fj+3d4LZve1OhKfaClixqb1g3PPK3K5jGVOfh
gYJSi2gJY06RFyj4M3A/CgXO5ufYCaeiHpywGR62x5AsPmHz9V4N1YUyxxD2upGheip3TrwOWL+q
Xuf2IEbqXWQRzPX0DxL7wRBDgq+iCggrTnBxSTU0ikux15W9ob1FTV0KR+EA3qeh0nq2UV5Q07Nw
1MlOd5SGiMknVsXKBRr8JUuHHJwMfYJTV1AWfRr3iUC+f6B7mnJn1XJT6MXyvRddNOID19/080tq
nN6kaU6vQyAZrQBDdcUX93Od3ElP3KOLoAAf9d++lqbG+ntPh7Ve9NrXua4G1E49s0K/sPjCBG9k
1yIoyqRG6Gq8PBlC1XnMn67//AZ9ZxO9v7YcSwOXqi9ifVdTOYWJIpkNq9SNPc6jBFfUXFoOf1SW
dLzIZA+mMoY8v0VxHChkvkv9Zkw9sSHfr/9mZ2fnub8/FZ8kh9JEPzj5Aalr7lEBooa8Q1QfLu9h
bQLWceEUPVJ0Ux2ISx6k9MMoRN/v/BZ/cxUo0irA1/3/CSWya5rNUlDwjipGxoYb4HuBL/wwd77m
EIIXuQsdcPFt+pWPDRtCqKxdJgiSihSTZcgwq/4K1tssLiU6yk+h98mfq72XUj8yncvFtSWUjfkT
ghtMbaCKB9rrUffwkfRhuSz2TjIs11HlQOYuT8jKPYI=
`protect end_protected
