-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AcSJQX9j9PcWc5jfPC4j2kzPbZGHPk8r8EaDCEielax8l5xKjz2T/yiDJC+2gUqTXGOrAFGpQCk9
NrIwZBQOBLVR9fLpODNA4P60SclUmS/5e/nNDQTXnVpx+c6j997VYqQUXrkzv667sdX4KwML/TXG
mi1dgvAenYns+Tq5ttuzkA/eUhAURGCktMYqrIscF8aeU4lsTRFfnXHw7bJ7ZKSgqBcLBepQcWb3
2YnPdNERiLwE+1R93fiYecTxCQVaZpJTQ5PsRJ4UcWjKr7+wSOJVcIK6Gy/Ay4bXlYROcUAGD6DQ
nuBoCg6wRGL+SPSmECxAiPlQwu/MAQC6tsF+iQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
VBK8+lT8IA7FBgW8Oron39+AdcSIo/GrornpXcZPMFhiU/HDrPLjc1DssJhRZVp0e7aAmoBnxrx4
sZ/wsDctYtH3F1v1fcQWF+eDVvlVin0kydw/Czz1DTDgf0nbVDgfv3KWSi7ETzvtvXylp/esaFTm
RT+QL2zOj1UbkUj8d2ugi9ncaWxrKI/Fweu3/zGIdZqj/h5rLvJ0Bggk+BZWLF6nP0445rt9ap79
6lqwAFwDMbSB8fu4VBUpRRq28qw2Nsa+LkAZxSLCCL7y7xGFAugq7n9ygO+5mUX/ea8eWi3g+1aT
ZYs3m/fx5glsk0yigf0jEVysWxwHNDc9gupx7wupqXFfefhedtTqRRVVQGqeSwHXM0NBaebs7vJN
fwyTKw6SzPvruEwyu1rs9CBQj7hLEhnmSQjbaz70/e9tAzaGBlTxXye/fUg6GR02Acd198Yv8zra
ki3JPJtC1161XoC7CgY/SsgkMeB8gHK9wxEb1acU2niSQ1QOMBqPLyKYD/LRPr6aDVm2tKgEpqtq
aX7ObS0OU/s+JNppak2PaRaoGetZu1VXtDZ353aapxGHIXSjH50W3uUvORYZf4ozHrdhkMTWy14R
UnlQKK0XbIS9wNZ8RKbyTUATH0TrefCI020zSddEr1QGeqOxhDMQceuzRpvFFoY1+1GPWG5t/1vu
ncU3TDS9QwaHPGYGBOCaJTHOgdjWjUZG6iS84m0HaDXyLYe+4eozFN+W2eA9i0S949FJBteQZWcI
Tzdfis1mMVoKJRPGcIUxkVlofFCKmOwkyAD9100WxY+44qtzIiA1jcTl5L1PcZP0e+xGDJucT1T1
s4mm411qtoQyl5kwXZSyvEmNcgNI5OsE+j0WXsxgf5Cm3/L8tk+AtWxvXPtcTMjuRZBfAKH2kqGm
MWT6aeQgY7j1WBZEbz0ded9v4qIZKSRt45obLnACJHP8f4cM3EIMe488aKXIoRdZi7/vVtjEnW4B
sPhLRbP1xsjobmjH3hsebh5wq1tpEGPwu6hcjmSMJV+n+6DAAu1ucJuWIig7EFLrGAkMQy1AJxK7
LMM6JljlggTj8vXR54F31ddW1+y3nJ81l9Y8qWiJP1SW6K8U5hEpZZ1+dAR2MdzSGuuL8K/pAMbY
MgrjWpROksAIs+WpWpG0lQ3uKFFUw4Ym0otZPqjyTRTiY/YssJ/CEVwnm+Xa2GwBepAl/bRmhFrP
7KSZNDU4oC/5PtlEhCCQdZMdEauJNFw9CSR5IdVkbLE5JY6SfU+422y7la7WYOmlB7P0MNIC6AGQ
NAVM0DzZx7YIfUUybYAFOG8HoLs90w/BR8X/2KBvJzUyIPSsi5jOQHDtqVTL5CbYqJG2AAHBovlR
XJDcWWTgCUPwAz7R3dbNGOVXZpCQrmFuIcMa1Rgjmy606G7a378XmOdisGnv0jSthINsYyePnHUA
NQMhQboEWeiky8lqNIavOjhTmANQqzaNzoY4B7wxckHKy0pFFtsb07hXWQiKeqfg2eTqym3Uvfje
4yuqWHl90iBX+50WhLdwJr8wfT/mpSa1GCgOxEC4Fg1btvtph2/pm9VLGgdJRqM8g2NaTpmQNC9r
xpl95Ig2PqwHuvg49qQSHyZEgLQOETByn7/BWGV6FmWSNfhaF22rn6n+ThsJutbBObe1F2GREhxi
3ITfJugm6DyLYfjZdguf8MHNymAkjNF/vH31K8godrmCYl007u4CE6x+bxIcYKSRytvyXhEhR6dq
VB8/gIXiarFCUbOh56TDXzO876t9SaKrBRPCPJg+9ZkuurehaezE1sJF4hcAj1eJlHpYlQoaxXR0
RgC38ux62SaT+fY3knXnNncR8sWB2FpO/qn9zcKuKz5c2+EhmdmR9LtroP84frJJ6OODvqKSzh15
WpfQbodkZsQyaHdGc3D47LCoEPCvm0pMHIXHBOXppWhUMOVH+GSzVfaUmlknGjpY+D2bdGecU8Uw
WALfaKQgrk+9Hwzb7+bGu+Wi+jB273Ozm7sm5CUiN/L7VL8yjmra54jcfKfQD85Mgo1k7SG0Bpas
V5U6W9uuBTvjtXdT9WQhkqb49LtO4TqFEcxsgaULwuclIzHJZHCuStZ9kLIahL7A+ZdZGImArIxa
E9MIvxs6XgCqpsQ40zoBlMtOLND6FUiIZLDQwK/K9WxuxwfxDfE0t1STa6O9nPRG+gYaRvab58a9
LtK07ew0da/+iDuEXm38dkzSM2X+adls2UxWncCxvbzE7+8hl1YkSE72nDNZ1ZbJgiX4pwV/qZ+S
7mU3FwK2HmKTGrS7HHAg4pqDSZN7TWGcGJ9A15zUvryxvVLaaIWqrRClN/WfPB8Do8s4XipI8ho2
nSSOFrgjeBuGQpyE9P5cfDo036qGZo3dPvcQ6i/q2H2C3mXo7lMOgjbTsn3cGdUset8R0mPLM1K6
T238xFPvim4IUtxwwaHTh6q7hh2vHWKQUfODp6juxdmX3j6VaozcaiGGXY4bdfAnRmrRjL1WF8h2
G7A1M5zJYJR1F+kNCV2360c1Ep6LUJkOvFG+dmpcWl6lk7GNfkaMTr3oJNtDZsnc59GJngjrBz8r
bd44uu5We5uZUrDh6VNa0D+3hFSvYMD4qqo9N288P9yhfUh+pFui9tjnKkB7DljVBT5f9sR8LUMF
XDSuu0Ak24ssq4BMOoyY5GyJAQkKXEzrLSdLrmmbvvly72IcWBboZ2hQ2JQjNl5u0lSATY/bNXpf
a9z2vDdfUlzqU8Ew+sq+ksAv0doePZ9BK4oTXss4y05rQO44GuXj5b1TkP5h0A1o1uzR1jRzowwc
V86Znx8b1UoocdsZ3sydAw+uiiZW51c/UJcimx1jQKJ0dfsSmf8G0iSzHzDcMhVvJWBMqgj3glQP
DS5h1/F5V7Uq+zPhUqF04Mp66Ul/FlS7kCYzICLdQLrDBiA+q1q1BZ++qSzBxM1hkNkxxRvCAmnY
XA5RDq5SyGHIMLyRSHsy3UWjQoGFuSB+YANCSdnpDfhWEHBe3LauwvaRr4Q8GIhCNIoVFBpIwegc
8eQ/YJd1MQIB8ZrHhf/KfcLd/JldB60iZ6e/5PAK5C7aD1FVVPSbYeOQJ6R9JtCJ+9xvB+oMP8/9
e9tsrmOq3EX9D7ROk6xn8ufzwv/CevQyRfq3Q11/+Kzmb9ou1uSmzATgQNlVzbbBFx5WzCi70hFp
gs+jUxsieH1FTgss13WXMb6sKNuFyOLkoJ5ceghQskJnMnNgeSQvkOy+bhVi4dmGJIZO2IIVqH6/
DAK//sQuwy7UhEnqdFSs0Sp0eEEhbjUAAfxLqr5Qp+OyzyZ1+1KuOe+0FRt4SF1SeFq292VWI+b9
IpAwywyOt1BDt16cYEqEhGF7hra8tU4zDCJ9gL7cwiwHsIy0ihQIghXKtDTv8Pn4sqnnAtdiZHHZ
uNKSfQFe3xkZX0ctnz18UKUjjc82AKeJCIDP5RoaCGFdHQL0GKnC+Ex4/lG0AeMnmUa4jeyFWpCb
wN1tZBGa2cgN4vb08oeP7nZVrXVqvhfCXcqr7g/HRzhy5ATZRlHYcAWcp+kWlRPvtEWiVNKYomKy
HIuQjs/WFaSxEcAOJLVPyDLBcR61bJYFk55+mKmlROg2QDU4IMO0BQ1B/DJPZv41+mdHRDxVRJmQ
CpokRUrnxtpCJkeZTkTp0wzvSLOICnrnYkPV3RKJY7vVgadBEwqD0PTJL2/OvfahdhOJpXviBjrm
+algfD4PhtpnyjgYzGUMuuVXy5BgbCCobtt+7tBcrE3ygkfUL4hY9MWA2O087kxVmSTp6etp4Mtw
kMgrk/g9HLi7KR9vgfUStsHuuN9PKzT31aUmyurq3PS69M8oQxfGSwXaukeB1s9SCWGFrLOJMk/6
cHl0arxYBi1ED/QChl10DphO32jRy1S4BkzrxgRgEnqVurcRjyyJxYb1UoAx8scLeJX8WL+wPZr/
IlWesAT794UpY2WvTiHTGb8SUTFWCepTbYFAUASPrs0MKyvFMuJtqpWKT6ISyZKRukOphQ59rssQ
2ReNZ9nRG5U+EGERSklkyZKqmGiCcPLEmfXEzbvFB5dYSpWm9vcGfMB0fBX0bHQBLI/rSkDyZaHd
mTEtxb7ZtjZsCdErx2fs/m37kgUqQVmZY2dxmVMyNwF6N0cUEoKIWl3KWaJuOWRBrPOaN/YtNERi
PBfbuaBIkeNq0EViJis+nvBcX8raZTeQ19ktK2S90o0wPYMZPxQox6vSxg6dbuIFTIgUdUtXtxlF
HdvabbbDVR7bUwfFmrz45eMXtbZATtnwGh4rfbYkaNj22KgNiFX6qoADvAkXjvaLxY7kdctvohU2
rwCgJNhAk73N2DJXl5IHmv/pVZA3vSoyJ2tdR6woh7cD61avZCxuaRD+HN/Evm9bD1lmYkMHKe4l
+5010tl2sWdQTcbLknv1ecEu1YgSSZ80mzuHAUM1RxSNiLvy3MNh2DsvpMq+7lJsbLg6+pSEZUC/
4TLmaMc3nUUSrjIXFo7RnFxFji9NoF5q2pqJ/VxZ6o0tmzqeb/LhbEPCbETEYBZP1LHQNg3gwdEq
/xH45U/I7t/B6+5al7ubkLgdyq+GKLMd/eSke5v1V50S5VdngZK0x9TfXGA/whvBm3ScMI2D3x3G
QDsSLtQQqIN9aZnaLEVOxpoOOAH1OQU2g7l4AqwE8h7gRJUn7D1xLul7gzVeB4+qEd8Iv681NFTE
cijUVgEEVpxwLRV3Z07G9WVr/rey+RBPjxYrqVu+pWoxfTZpQf0fj1aGmVDZKBqTXBWI94ns4u2e
BTf7RpKseAlGaxPTjuM0xqtBMx1FboLIhYaz0xoumoW1vo3NKuScfzhiTm5wHU1fpdjygttj7n38
d9xHqEYfZEhJTqTr/P44ELY8RGqmpIgXO3ZZBSQ/BbArK0XXdzSasODXgdqE59gBqFvgcxO13/ck
jEbkeELCdK6Y++LmuuhZ88Ti0MuRD3jRcQMf4jRBoW++CHzW7TIf+38r9oUxx0m9d26uhqllyPKx
NA32j8IvIT2ynh2nQgPVyd6X1PdhmcEL9YuIf5JT522G9ExieMabHuJPLwjL4A7m1IBIrRnWSWZE
GB862KMvfRjL3pbwYkm0A4WU2FHu8wH2/I9QJmWgpp1BlG2AurV9zOUbKMWWtjch950Uc/lDR6+f
NzKzGMtebC93YzX4/XJZ9e4czHC1BWlGDRAR7n9Vsp+VoQwnii89RnO/8KG9SN2TST/WLwk4T3WC
5cklDjrABFP2vxUFFo/VVNzgXxLMTt7ll/fgOsnM61njajA7BCnd1HumMkaEDQj/am5GObsP7J3H
HbXX5nVQ58WAUMksjjPy0lM0WAU2+gtxz0dw6yOzQk1bu0x+KQZpa9pRGzf8gTcIkp/43AuTkkDb
I3ay061CLJGqHpnB8LHwP9N7are/QQOaEU6PjfjsRmECB1Gjk6tdpjUrShCWMhJmUeV0PH6Klzg7
t5UpO69W7H0I78B4ZdxPVaJ6rr533pXsuUe2U1oZU4sJAulf8zdblRB0uGlo0Sh0xhOyWwX30LNc
5VB9tU5zM3g7PAW0esUB6tVbPPAUHuH6OJP8KgzNUt+zgzwdsFdAA4UEndHy+ueDnGhqLa0fOvVL
VBgyNiZBahvaLZ+d4RviQoEp+DHjnovT/Kx860R4Jf69qdArqt3QKFyO5V/uVtbL7t0l5ByXCOOG
L2hULUSltozkhyJFWcGh4344lsmiY3AWSHLRhZ5yEcjl6pcctHQrZCIcE9oC5dIlQeSugr7fivJ4
ZrKHEO8Md3KhxYrjb7BwL1uygPx4MJzs8oNyeRDKM4l5vqhFw7HqiOW2W9WHDASqEzjr0ZakQMAa
FhestmVuTyLNwY3tg53C+WGQk6CMbDzEZdA4H1hI4G85FDTnnp+rjTdiuD2iy2FgtjV4ef/w6cx6
YqL+njYRKykRLiZzZxILwUSz0JgjcefdFWa/yhQdK/Bn3aXME4ADZxxoF5EUmZatTVdREpHwBI/G
1KziyHZ1b7ODstSZ85jq5sQoRY24Z/UgD5KZL8jWXowpPVY5sSwSQDZEhrK/bXQGIY4D9t9ZCZ2i
3O+i0bPF7cFJpQKDutJFJo9eSFy7aLtPy0lfaUQWdy7nP9Rtxf3in9Nui5b75NDFKosvFn0Db3ve
eBQvL1vE0BFNv+94JV0NjCJShjwH1D1DITQzXn4eFMFn8rmgS4EvBKI/hkiuFwfXdxf5nSOHALwt
v94Rm1vDpJ0OuWKr13tkcO1m+pAI7GWNTHYAbm5igPUAcyLoBh27R+iiQDhPZInHJkmA7J/PEW0t
HOtc91ahCGMcnhhP/0HQyh6RqP2aO0vquqkoIX3kjdsyPoWS5+KxBvh1SO3pY3UzXXs69tG26+Ap
6qZ79l4++zS1ZJEamZX0Ioof5poEZRRrvf7OIGXTMOSaA9ih4f5FNMs5RTywPcQ8wb7oA6wEL87s
NFJmoJQTniH+Bn+tCWu5o71rDbJyohmr0DUN6olQXSu9nkmbGq4hIqmt+qNj0ffch/3USIfhScmK
3FiUsizCmpTM4MdcC8zZt7Y45X5UMQZLP2cyV2fsigv7m9Aq9+TpXobf5ri6bM6Bmsy8DHpz/xgX
tF+HtaSO44z90rzIZmI/mhnJ1Gf4cfR67Kmqmm8I6+vo4h1UwOL0bETfTeJOEEM4S4x/xN5jWEUk
aqfbSw28LqoTkg3o59DqmZyEyoiTgEoOv0WHQVUpgVIJDzfoC20/IhD3h2LMqT+WY4hPgDJnvdGl
vCLVcSZZQsqe0ba6Z8s//stThbS1yBYwo2NWMM2cTJ2hjb5jsDuOqZZqK3sHHfWomFDUHGjve/NG
Jvw4yHpJ1cKMKUmieTUrNNmEkgnerTyVS7D9Ch5q0PNE8kSDbl0cd9Ka7jvRJnyKygIpb30/Z2HO
MU4m+YRn+IndglQw/T1YndYxOBZNLdw2QfKV6RnLKzDmiiLBJ0XtJXwNSJyYpjRPzWtn1YbyonkL
Fr5fQJYeyvf+S+yQ9bQADGUaywKX7TfPsVv/p1Z/JlSvmF9InTHoxzWB8YaGhPC7zitsrXz5C7NL
fN2zsgye5ONJJg0/9xxu10vyW2LbcEs7OlkFl2sPhj53HEepDAZe5iLEWMLDvCXGg7fGwF/IhsIj
612gi5V9Lm6i7bxBOjUrXAFqX1KxcGg7/Upl9AFIs7gc8z3QfXVEla2U4sUI86/WhH3d6inRquHA
hvZj//EEE1TuLTttuHelK6hxkNZhc9WWge8vf6rbIfYR9QWVo3I1zM9drPW3JJ/UFX4hsUp0fF9O
h6fZoXZbgxg0+FpJfvy8wEbMfa2YRClFtbNRorND8U5n066sBAI7KBzDB2RwHWzpw5c1Oa0zYh2E
UGcpR7pbvgJ48x2wIZRT8dggMtTiOVTB/OfZgG+0/F4oD9ZRoXiRktDv0EeYglwrnxw7i1dxg222
e2ymTSr2mlwaNsSbzpQSaWps8SrcBOo476NtOCUC0qFZ0Xq92iGkz4+q2p0u8daaO9FqdvRKy4ed
Z4IMRKXBa/XJuyexrE1yW+Nxh23SDH8MGqFqmRIa1UiDaRF0X0GCo3TPlr1dFUaaTyxot1xb/GGW
Kpj9Sl9+e9xCt6YnGtMVUiZ05pJChiSOmJou+w20W+6zwLwgZeCu0XxqdJ3Si2cbL9+GfV5zBEpU
SSCl2dTgZJQrcNOT4zOSc/KyFIrfD/4R5l51Hk3MPkN8lHhYXZfiaTkKKDiswtUbAl1pWPDn/k/Z
9/49pLe42CyOI4sQlUg8DlH6UHbMkLBfEoI9TFTdQ2MdeP4b7wG1cRulkHmTAFr9rvkeDRaQWozh
qpTr2d/iMqCUGpED7jq7Qn9aqp1ptgP5kLWHzmxL7p4VuPFa/5MuPnL91lRA6/2Bt6vwCH45hn1Q
j/+fhCjfiCJUls3ml/azmQsWQNAddYLBFFi2QXVJWZ1v3/RcMFxbyBrh5Um9xoKQuSExcxJg6/oR
UHz1mrCGf+qH6gV0XqP1s+dvsP3+AMoRaovXh+Z/9eyO+x1O6DiFF665V9wKFyjAyFiqqRCzH7hP
6KS270MvT9i9ew9SDvoNPrmLdywbjEXEw3Gk13Miy0Hqgl8DHptZNSAiBXOO2DqbUx8udnkaPuHC
LBKbMmojhvfJhmdaGlWKPggNshc1FQB3Tbcf0lOVZsjcrocTt7OXGz5TLoApm/hOg9HpUwauzmA1
U3OBja0xcg095kuKofxV1aEqiooQ63vUKfTCwR+3RWVYL8OMoWvwNrR6FoiI5wZq6xHm7zPojO8g
eCmnFiN4IE6y8Jzx98Segkf15LGWfsdgtqBcTSp9+umIy73lxeIvEp7Ea1KirKX/AKpvDY6vi2qT
7KZ+6523Dbg5hGSru8uF2Q6nu9vkYfxUbkRtXrO36aP7MYuCFFMvehqXgNiv+V4TYMyMJSM0NI9L
Q56tB8EDc5tO+khkV+49clobeRTt0GTpujDUcOWq6XYw+Bzz/Qs2uS51YTtdBTpkO7FjcekRMFFj
vXOVUcEUTvunbmrnlN537xZFQoI9tpYLpkXsug4oc7bgY/iqZphlT1oARMi8NaJAjcMpJhPuwgbl
9UMddiM6BhJlHbpei83tVdaqf0zzOLrE8gDk+7IAP66jszwEzYST2QKawOhTEnkoLsLfe6MJa26b
qacJraxlh76quVrceTGfseFtmhEHttdmIGQWI6mIbCmDGP4kSMKHOivQe7kYNIPvFMJzW5JIGxho
hsmijNtsXCzymH1e/wVlAi2gDcBWK5RKjb2AEDdC0QZrxUSe8lX+whbXVHO4s6G/5mJ3Fu7Tou4z
yOWeRhBb+nAI2LpR/fEQMn9cyNNevKVCTF9c6DDmvWftLuAdYPEkwl0+Ek9g0LugHH/fdvRdC0wr
XXe6cG8LAIEb0CBpBt94K6C66YVRHKRbNXZ5jyw7lWCbWWOo2EuVspwCSwVibx6R3m3eZPr6bOWX
ej1XN2c9PYAfsC24n7XhtvTmLYbr5yCnmFrXzWbeYVFJpgUsHaRVQ+e290cadecGEwrLPlCzVBxH
R0WiRUgyaJW3snOmgmldeLqyfxric3kd0Fw1kZ43x6E+JMdHNOVY8cIBFTuDSPtiUKR6FRIXgI/f
NeyqVgIY81KpaKpBlzLYau4VUqI24ow9XDdr0DMmOWZVYhpw5ayI8ecJgTrePGiHnxgC6z9mXIY+
wORfoALWj3xQYNjrPekVDsA4KtmVI9neUVRVs6smzOizGXtShQaTr7Wgw9sBUO9s/Na9e+HEg571
Opm/HvGhyNJcJJlBP2FPKr9bqYW/O9f5Pb0d2V1Uq1oFJTzj3wGMd6QrrTcTdpnlUvFnzi844Ezx
Z6JtF3AQZ5dYqBTOoER7CHKM/EFEFt4T1yGd8KQUM4FTBLPPh7jbrcjsfjqoK3jCXLTO/xJMfuuk
XgB3lI0T8b9ADL5pesO9LZS3X75TPYyyeDfxPjLdpEdzWo+hJSLtkErhc2nxCgBdNcYfUYt7W3Lt
w84dAHi4aetPWG6wYn4P2fm3PV2xlsCGYddDt/HgAoidxQfO/4M70Jm9AiLsmX9HG/qOQHH7xtRp
JEBX1fNmpbGMkYVadkwi60W9vbijTD7coFU9iO9cLPv1R8lkopoGCHZs4tWyaAx/OcalI+8tzTJk
jgNIMtaLVgUwB+CppaHAxpY20/Cr80lL8MHlnaqxZx3xRXktbRXvKkG4U5vJL5Cs8Ov+ERGh0MoF
7Yuq3Hb+oRfCiSIzY/yzFQSUJHMM+RL6uw/17ENYE7z4xaxRpMk+Xm636DhGA+NkxZ50EMc4wQYq
l1fdaOH+dxMbBGLZsJvbpgHIVgmxNO78HaE55BSdDvjimTmm89A6FBapJ1Nqd4yM19RhfKLGKe24
lczRYug8aX6O+yGytDKhQ6Qt/F5/Kj9GxlR4HdtKSqv6/y5F5hqi4vpIKEdq+ghkdTWKnMFckby0
ouAr+KfOzXNI2ms/k7Mf05Djx4eQ2Hvz1N+9YFyKLltX116VvOBOj6mkeVWdxOWA+/J96H/8LGWJ
fa/9DuwgNFCrmdGOcNSYzJqkH+WSeehEDhCVkjZTSDvWp64YIHu2tMW8G8vZBfSRXcULTwuZ+EWZ
p20TcvYw4M61ef38JyCpvMAUO3xh0WcKLGDqi42ZNaWO5dv7xcTqXXIda35avhZSjCbn+P/ZpDKi
5AWUfINPtf0KrFdk40Vz0o02x9AGbxYMy2kklrFXNQaiqL+SYPp219n3+0TT2GFiW3kbT3+yqlY4
/Wmqw0gXzT2p1nB6JwYlP8kOE8NK68ufVO7j0ryo+E+EBUPZvXl7whgQ96JJMQhlG4+xYGzHR7zx
6kNhoOXvGNi2WZqOCN8iiagFgCwaDnwA3wkEaHh8eEDbV+5IyIwI6g4/tadJ2lVRkra78dzYoyg7
lu49Ze96BWgR8cETzbOg15m1L8d8Gom6FNHPO4vW0bvmJ34C+WpU7zUC39TOVG6dQZTJJDzZJFx7
am8hZAdx99naOhwPkdsugv1q0SVn1D2UMXWLB9RjXRMhE+82zXX9UKj3nNysJRO73zoE03so/bmC
hSOct5BiLsuTPHvA8PK7MKsVmhjCyH0zKu/PfT8jeyvX8k0Qr+5rmY9IAaF7is42y1laxb935BA2
tmghybUUNE+GZbFJsfCPAvw3OJfLGiicA9hdj82CTjnCOaHhpLTMmJRfMw5sKrK1JuvK5MfK7YdF
oR+/zhhGod+1z2PtImzkJmIuTZ5mv05EsEi+ppQDyCzJaCBVeaH7235cf+de227skWvdC+SGu2O4
zKTcCZ2XoRQ1yIDeMam2n/O25D97cPg46QM1jxlRx1zjhavEd1dNrHh/qbq8SfCe+v7kkR95PaQP
Qtp5AB8zuVbEm8uemi3j70BidyTT4URZFW6cby21fS/UHwoloDtD/O65X6xFAfBzLhQOPT68py/I
Vb9d/p7G5rxFtBL10bS+6NB44gkdhAGx4DAwKN2pnEDUMBoz98n5Ur0LzwZIInc7WpUUtjFMJNkD
YEMoSH9mGcFUA3Efhb1DoFtwCeBSD7e63uZzXdWwyT4J6R7I+qxtvS/wewCUi9Pf9Im6mvNUeHFQ
tRFAcEpAjxTrQtSr3hpDDt+9Xc6lF5wQr9A5rMrn5MGIfJeKqkWU02HlfESkPKhcMacfhofrbxBK
LbioUuAvCnP0qP7tBFp49mPs/UKJYcsWmedFozcLSgHs5PEtW2oEi9/PoqAVSQqWwSRvseE+N9Qh
DlkW843KwmbRsj1+wS6K0BvAtz3jbk36NRq+hjw5MfIb16Q+ZO28jOMHmgWVZ8M3YpiluF32ba2F
vLPxg0TvsqHVWIbWsC6Ic47VQ1dRh2LuvTfJccB/kmKIVckTDfRz8qWuD5yPv8XBgmv6GrVCK2jZ
LoiVUzyCNy83OBMVj6zZc7inE1hk4DT/Prul0xtM2pX5dhEGtYxTh+RWxS6EEb0juvBYJzJCyQFl
gyv3nN5Us9iaT4CBWD+FExee64OnZkHDsJmjW08Ob2kA33Zcvyc04QCvOZCUzRFlHVVBqMJMBoVS
e0OHQ7qSlwLJvFBiyNxpWruiNg9DjsWQ6v2+BH5h358MuCa6RY8cJJCWOWOWvYsezRBxxmS6W3MW
hOUA87Gohi6vw1WQ9SuQLbXkp1WoQN9RH7F0dMpkcZE9QafVdBj2uXQEK9dv3jRzta+ffnmZQg+B
vTYQKbaqPrWLVeeAlcYWF+HQxdGcbnRomV0MBz4pAllrv8YcdcRTHj1llahzC+zRJU9H8+8mbUqM
enE7FRdzqLJsZexxemFqbFhAjXxWciGjU8euINGEzri0GKTMIZxzTjsxomvVHtQD9lvv0GkCwl+K
YHF97Uakcmk5b93/pxFYtP0551YLkHe7hmfY5zmovrANUzgIV63fzRcwMsz32cWAxjlN6fMVvJkk
XiP7EhVvICmuaqa6A99iG4kMJJnkEc31zsBIzwEK4rBq8etevbVVAVkhs899wWQHx/w8uRB9hUeo
1NbcVDoXe/RvAa8e4vewUQLIJrbrvAd7cC9uxZdWXtOAwVfGLv4rb1O41nwxVwB8txuT9featdrc
l4SeEtO2NQ28YrlcLkUXUTF0Eay1Dc+ptHlGs1YhtQ2HXGoGSPMrj+Yg/qXgB3jKoErny0yh1Nb5
pAPrv61+lGXURokOolHrbcWyo5bFy4oHZnj7PtRoISnBjgCWQiTe7GN8a3zAuTxy0AfhwtpleN1w
pkpu3XtCUiWNBk2d3Ot2GHX08D15T48VIM1mj95dwVPyUe9hriQ6U7HJxEseqW5+i/kR1esjFfDN
em+lXW5HpGMbFSik3ON3JPLXgHlbXSfuSPy+dDCBwAhhUFYC9KD3Z1s+MT2G8Gf5V3i4oqPfWmXY
5NpYYqVhgyfWxLz0+3Bt/mhcgGwmp7MnHEfuVagxg+IuEx/U3h3/1FOJvvUbbDWdSnik9FFnZi6S
kVwWzIvRkKgn2Uyw6C5bLSjYG2Ndo1um78SnmlhSQCCslcoRgre5tuj9XA8D6gd1Bd+W7DOe1dZH
g1e0QUh48znF9UMhtfP5wp2aRtrCZmlLno4r3UzR4eQiG7pvi3+bOjfmyiJevqP/bXJhPftOCBBe
jGSZPBPKr+cJenoGTmTCw3Z2bLJb73aHbQ7BjwxnOfBCLaGORWZDwpQ8TegiEKPp0KcDP+iOSn8L
/n+Oopol+J9AUk02eo0TKt13A/zrUn808EPKfS+kBIrwaMZbig4Nu5+WCkSz1UOnRsIMGqWKWvQO
1OuSuN3iEsonMXlM1FzLyPyHuZ33uP4hSbwBaEhPefKh0J5KM2n1AIAbJxmCg98YtFTks35zZEc0
TbUc/Jw3dtCika8H/tmbi/YWjv8PHyU576pJLSxD4EFi8ihkRA1bZafqpbEedCBz+Xk70G//X7hD
UBHgf6pAY7YQOr3RkZ9Q9MEUMlvMfiNC3XQecAxBawy/+bKy1L3ggvizqeFwpfpO5kd5AU6y39o7
K5qbjvPhFgsXjdH7PsTjupYICKIK2D4QqSEtPz0SHsZDLarQUyVIsjDDM8ELKMw6AXk6AFDrBSr5
bA1NZR4fdIudwa+bPR7ZSGLLTY2xd+Hmr88sY6qGo9zzCWVUyxRJe4pwpWma8/3oZBkc3Ab/UPaY
EfAKPJguhpJarAh9WIHp+WFKGAXFI/ncsyhvPA5idaBxwHq+cp8367YBuLYhJDi7ZBuEtRHAp9wd
tT2fuMcUJcXwT+sB6OKAZEnBMYQHbSI1aGCtlFwOIU7cnF4e0V7yksWLiDLt48vGIHT1hVncafak
maqCNcQ92JwmX2b47QBRBCD9mNScOMggGVNx767GLGJGviH2yTzfKCH+sxzCXm3d0XI3AOHtJU+i
aNN+Exfswl40yrOxQBPjJTjiVaEPhUCqH0naPbrSi4DPigD3e1bi5cW3BYmQ1CGOymqbqXzUxEvo
94nMUYlztjhU0bjvBLJwOAGuZJXN2XqhD43FwDyMUaOsKZqqNdx0gwCLWChL3Yzhw55Uam8ZSJXm
klKLXKEXMldWTP2xYPvqlKYluQv1UeIIxXZJkv+WJDVkDhzL5jlTW2ciP/805kTJqJJll2QIqv75
kCJiPKAxhSsA8P0stF8NUk9bJTQx6nIiwEs1vS7RR3luHk3n+tRudKNPNH2/Le3xyRFeFMvnLfSD
TgeHJzBboyKurTvXvksqUZOsI8XiFSJp1gMEz41Kl7szLYDjEvHnDZsXBLO55lg9ZnlZpxbNefOt
hgKKmdTx2oy72PlJXmC5QLZrUH6IbBPTZcly0CDOSi+YSlxqqANO1vaxrcYeIDDuFSKIhZPAIrjt
vWwoX9xbjV+qsP+Sgu0bsw5gPh29ee8ZfJNbUZ/387WasyT54H5RXwJV6MfIH4IxAcSBgEIszkzL
lijIX3ntcTsG42QRE60BCzY4h/A2cKw3VJdTXhvB12h1uOvUes6z7NiUV7kR9ko4jfrBW40U1A/y
5x729EZunhKBdNc+UBoq+n/xgslFNaEOg2phsL9ROYuuE1SvXMWx+fhLu9XHq7+w6QYgYJfwe47+
EYu8kT29ehKiZbhRHDmC30Mo/n/0LdsRq67RXdvEEpe5Tb4bQqOouS5xNcZspsRQX3eYV09m79D0
eV52/feOEHP2jr+ewWNIsRGj0M2RlWIL3CdVLIgUTGQBiiz7nZYb9iofUu/nIJtA4VnGHybbzoSi
IIKei7KfYHeYFO43j5l+vOq5VpDAwFoytipmGwDIE60ODhCXP0e98T6JfBuomnGd/IjsWKLkZWv4
g4Rul9wJ/U2XIBD+xYd30g3RS1zufSc8m32TFFA83ZG5F/v9/vPt+ouCH+oUIiQeeIHdORd9c75G
U1TVPKoNB/DZ1nyjlvZ49+5GLzUlr9Ce2taYepwr/VpP1OpK1ejzv4szSlxL4MlZvJrjnVIFsJkt
cRRbNg8fWKEj468ky5t72RQnDgIoJwhMNev5nCB8PN9Ac8N8Th2tVtex2VjPCsfhMg0A1YDR3ecR
T9v54grz67WKJaIUei+my3NpY/ZfpVmpA3U98d1ZN/815BK2dPU2pUYiQ4FsPf/hij/fh4Cv+Erq
QY7rQE+9tvmnu3qlOu6OSfqjX2Wkcoqx7rfNYekwTntb66Sas88IvbfDm1cjP9+zDLT9OI+jWZnv
tjeX8ZPQTmlRk4rsO+H44KWJk/AP7uynyYYPz6MPb2gh4wUh//uXqYUURZig/xdOJeKCTwYz/H4e
KUpEa9FCdF0Zm4OQyCHdm14bP6Ay/ipBsIw0Y7oAnBEWBVBqyXeSUmjsG63NPewQUUQmcNmUy9z2
MSbgQqrJnBPmww5qlxKYblRrbp91YX1zQs6cker2X+Ki2MeBHmHKdED7x+0om+i0hCc6UjjRfouy
5/2MjXa0hf4luiXYJIQHJ4dRigsb09ES4sJY9CDUajwqW/H7fSuxs0hMss6yBU0tHsGi3OvbE/OT
2Bo1AqaIn/kBkMjoylOjZWG70tODU1us6HInD4+SMqy5yCq2gGG2/TRpXlcj61hO23rhhoQ5PvBH
tyXV+zszYB88bvPyStZJfNDt5ukwvQW+uaWg2BH8nLSVNXJ3QebyfDPJkAIDhyxgd7HOCy6Q5Wkv
d8oo+n+5mjovw6dUV5w8Of34gMMa5RiK7XWl0YM/8Ym9hHXtexQW88Shiy6VCOQmMRN3NjmHuuUW
8EOzN/EuNLZ9YL6SP2/6VUI/kOO4fLS0HSAl8qFF68TUWdCVZptqAapIM/MEIWijvvFI3JXwMudf
wzCOZDN/t6yypJAHdsmzRpHJoY+OJN7H1d5avc8Gthn9Ej7tj6loFLm2IdTaldJkiKy46azaFmZK
bGew7sHNEOJzghUEiSJu0D8rrsynqg+Px6bb/vok5qD/JXm24XN61TCWW9efsCX2PXx+1/S/JCOI
PIHR0GYFgpj9jWThUX97BCT+kyrzUxXWVVCsDSM/zZTEgPA/dyntzOkRTgSN6FvboGdoNiL5Jfa3
WsiDQuyCR6ItgtLgKzZLWL7bFyfUerJGUm/RfKKmAKkfdwmdUzUTLUZHp+aKZfVedoDnp1nZ+Lyr
QMtay5U0o64XOBS29REdYHFN/wt1+jZF8TYIaYjIG1beGQALwMzU9twi0Xtsxh8uv8JipO96/6gx
HTaOBD8IiKLSbLwQYaxtAmRdh4oqIA3pxEPBK+GHQRLzWjxQCAki4KJ9Kswxc7F2BTID35h9w00p
Rznf3Y8pu1oSDS5wO0oRsGTyGd5Afa2l1RwEMJ8EEJpFfU82fdu/JWCEVFyLf/IF+/8JvE+0WFe/
m7A6IYz0rT+J10x9jqq3Fibp4yA7lsEfWNp8UaGu3otWOMGFBDVLfIiqPP27OTQAphgCzbYhOdGX
0sMlKR2N32RbGOsPYAF9zQilYW9poYNqI8jbSQ+THbGfI3Ykcp0NyH5QcQRo3h05Pby52orhekVh
t+sim2ysJKm/EQRxC0M4H+L/089vPthuhm5jddMIXhc+MjB1hVFTEe7J8Io7FVZuOyjxF0tBAvRD
eQrqQgJZml49+dAiZSN+tpA28EDHQaQA/i48QbaLZ1kvUYLmwQVRr3Vaa5yoTo65mi14V3qBkUaa
9jYHH3Imk7SBOGNOHGYW66BjvJDOl4T/RdHcFqRfPw0kWOgFQsoFfYAGjA7ErV2cQqvz5WL6tVWL
lK3jjUA3e/Qnpk9C7kh9JPl6oHedi2txAXrKLnHXDhzWtl3ceZpA9weel/0wDr2nNapSNB5byhGH
DcA1nA3MYjuq6tuaqI9cU6AXskTyPMBii5TF6FliWzvrzIytJcarKg3bfhmiqtTpJb4I6icuelYi
P4+w0wBBf0XPQBBClbwcjsYDvihJOMI1b7SyZfVZBUjB/UJ0QHHxPY43FDSJNvteoMq2bPNxY3dK
8GZcz+EV1RLua0B3bPufnzNiqxU5Gf/KLTBpLDJFtocNtJOQXicFi5X9bHrhZ52Wy22RxukvcFrs
p/8wEt3Ne8dr+lGfDTVcaobF9MTD0WtB4LWWcgcev/HG3H1fv5OBsD6L9Qu0ykPn4kP6p0dBuSCD
EwieuWqcHnu8B2SE2SBF0w78blJhw6jRdvVYFI4MDJanbtObgh/qrwASPjWGM2fwXj+N9lygLHpj
Yy6bWjnUeaxZJaqKl1Y1z34inPuXEZu98gz3J434ouPlxN0lDcNomdVhZ36MyJO0+uL9kEC2uk2D
q6gaaz2atraE30yefN4dRBS6XNrq8855M7Z6SJvgM167IiziHpQn9U6gFfUBgUT+nYFTH0kJTCws
58Z31XA618TQ9aC7dwwOrxq+V8pQ/47c/6CBlnLp8Xw0jSyTzKKFuNe5XyyUSiqDgkfGAMDrumUL
UipgUT2/xFJYQf+XArVngU4P7pepK8VaIiu2V3MEL5l0hwAHgvcEv+aNCL5L3gtNDgZYQDVhSsKf
MRy80epXT9is8m7Q92XLsq7iPkH2k+U1tSzNPEx/cWLUUel4KOTPnpLlw8jpoccmx7XBe4oVFEhW
fPt57xy/8Mu0mZffnw1idfSqBkjX9C2FuQiXVLAif6nui3aYAsIj1l8Wy74REYeoPMpgxLxYd9Bf
x83uSIfEX8NTPuTNZLvH0i6kz8zuRoFZsIOZVpd8Lt/Ou9Xt76J+8bquI8GH9wZxJtVTGhMrVlPz
0Yy64qPm6YnAV0WrugF1dsbPI0c45EUKPXcvhNLoftroaQLsWfMJwqExcRRnWgmLs+/NXnPuxAbH
lHjd0pDgZ0dL/dQ3Uz1cC6IajJWngAW5b6xMa1TgSk21+qXZfmimW6FDTDjk0IgFwtPYO00Qfl63
hgOR7ETDXtjQpMpzGBJw1NBLv6g1eb8zum/d5DQy2zZzkQRj7RQyx6jp4bMNIt0trR/j3ixI5OtB
TRBXq8lHNJu031bg/8N1WjWxySqQWJbT6ydeHmK+gH6PHSGObs8b3XJN5/O6+aj9Qshv6W6iVRt9
ga8f7J1Cmko5JQ53Rd/rar+RDglCWt7yiiDGi7InJzOCs85/6zb0cgdWZBVCzBZkRG/+jhXztyvp
8Xi+DMqlSySPoyGn0Fpv9xVxi0cjHODwIrWk43WouKzbnZUEITdSbm2v1pNdyORTh4fa7kwa8Gba
rLrUi23/tdLwgCvxsOhGt/M0Zc/FDhZ36QcGsnfKLehgIjRhta06lldSMumrM7+WqTVQSHGfhr2c
rhFmrX7LGAoBgzE8IxjK44zR8XBEmCZx7BFdkPlAD0GhPs/kYO1b9nk3/jRWCVsf+HMpFnZ2xhoZ
YK5PVle2N5YpRORl8qPEB0HHLUyRF56IJ98IBWmlVEnPysuf5nqFAKrPsT3SBGewFnuxrayJpDnm
l0Ebl/Y4APg+u1qladQS9hsqE9OJsRhtwhBbDpAS0d1nDhkOvlKrWUpXaEOcImXkXCtFEABq3ZWV
wQETuLjAQyX6y+VmjlveNQhXqPNGyKHv8l9OYugNyOYV3LFQ162LFMmvmJ9cjrpwb8066mfFtE69
mDYRqyHtWtxDq8ztgexyM6Z2oGR0B66pr2T4KuHR8yBZu6+bBoxpT5Ex4i76GAasWcWM58oqZLhX
qWCu0NgnvDOord8c2Zhgj8hcG1oP+OGYjLoh36ftfbFqvD4ibjAmNA2ECC1AOJ4c81fRJcmdAx3P
3svFwUkzQQsnUYl2rbelg92fELDhtjPMsvq+KbbLGOl0vwY64HL2XQNNOb7ydSRhbGf5bTne15WL
MhVeei1z9u1lW/GQK2Qw0YQdo62yTJ3c7GlrT/41SK/AZQcl0c9TAA0NUyZfTAUtqr+scTE/7AUV
oEmGXlrUpgm4/JOqN/t4jIv2MmhIyyy43dBVN4H9eXT23n/Tmo3ffQjFHnR5/05URmLUUwgJANSp
w46vpyTkeHFauhjP3vv/KlhgBMSkonhbTGsYRpNUf6NTxzVw8B0EowJklSgrRoS/Foej7aOsfVG0
1ZvR4gySSyMYbKOv93CdAaYqdKCXZjMuY+NQ8a/0CDhdLxAUkM20dwaBpkBFqErrVtyPK3aiTx7K
ZsKwIkKv+qCv40ph3/kxo+swcDsNwUuKwSoZkKjNhH0F8/nKfIyZh9Txy0+09Cerl2uXcBAb4taW
X1vbE7Ut2nUIpEPVK+NXJTgNXw6WBKAR0PbXN2PD1v6sNjksXHvaWIY59OnKvlnopgZ5rNFozqfo
V8w9vr0NGH2i6xTblqcznRirPqWamxuPqTc8fp7k4r/D0XtTPxF3ThVvq4jZq0+8XYs9SvfAgE4S
jUhnHLQOFTbrmm5ncn1XRXAeTLfyDDdwD+N2Nu+A3NnyDbEPtlDlGAsE6pWGYDpYPdGrdJ2HhUTr
oif76p/nSbyDeOxpntArmh2lrpbKheOxmgtpAlHM+oHlVEUcocXjSQGiTOLfjI8nFZtxlce8e3K0
Ip7w+oSWNI6bJbhv5RAcQErp3wyBrd8xp0gM6+HYkhDGXhSdEiS9GyTqP3KNgmt3KCg0LWutZXPU
12Fh9dEFa6XSUQucBwhKQAJhCXyoIDmZsj0is7/S1vFd//BFTahA4bl1kHKoVFrdmn3uIuD5tbtN
My9QbMIjH7IMu4kD40PZ2uFWpwRSMjRRxvJsTxFSgqreq1D30RJ0n53B2bQb3ynw5G5IjH8LyRNP
m/6G3rh37glP64YAqrH6OwTk/B+iS6TH76NfFNpetQmqy0WzpC9jsSaZYJAcU2aOoofR7ojKYcTs
28V9vXdnzdkz2G3/TWacTCfXvUOAEQdH6OoBBI/rcamQ8QjpbhOe1/i/NpopIjDc0DdE4KfyvPhv
y6WGgwOcmEjK9AS+YJh7qfi9e9x/PnmEfjBXIKBEEyHElFJyXTRLcU5PlBhFtxbOW78JtB0K/cQo
/YEvwMyLFxrCO94Oz87X07gtkMW+ZizDHZcxMcQD5g8UowZE2yIYrEbVFpul33MSqtPvF/z4ErwM
MBG8qJ18WbpJKey0FMVVlE0Kx1KgQJawV54I65ViP5SqwhUdd+/GVZOkGq96LhT35rT33oQahmR4
FdIn53ZIwD0ZvfQwoGB2mqVzrcHHahArOBB/Bdt31tchRDc93DYZdxPAud9oUchFCapEBtphM2Ti
GfnNLptto8Fd1Z1czBsHabBQfsb0jhn7FUWljYs0pJgDTQUf3dpQzTK4cIhNfYLZXv02iJ8U9lPZ
yLCk53wUKEZsSmwRHr+RJdMl9SJ3gjiPu9cFyiJtfgZJmRXopWAt8oGAMvoDP/IbfQzo4jvVDvLY
dfUazF8dkwhzr7eU7B2AJJr/7BIZgWwrocvv81uXJmzJOU3JS0kDg/6UvibG8c2Cvm+LTYrN8rEC
SpZW34XwockgNGfUV4yNVyVr1wR0lLt6ehwYM/qJwF2XCKHHSTvxgbu06BPYVIJnLvCngC/Ro6qX
EfMhqhbZ9KrUi1xn4IUYOuq5gX0bbVkhNXin5X6ImmhY2b/kNBx/rsH90sEcQnzgje3QhDgSrJMH
Yhkpf07ip6ilfhYelAH2cYVMVpcMFSq5AuK7SWhL/WzMwBxKEDnP8MKm+Ic/Dv6Ro2NRB32LW0rw
2Y8OQ3nwZCLskOQSFF0oZJ/PI8H3RlAOGJfdcaLXofEkYm0sHRRAqNWlNI/iQH54SJVGoVDP835Q
6gAIMO8z5mFlorsmNPCh1flAQhVAXKoAcuh+VBpY60ob5eAbP8L2u/Gtdxon+vQmkmwcQyPQO5MI
SCWXgeYkVkri56YfxwDcZgXxWZeo4S+bZmi14/JvLjOCKlMQq8vv8HFCcggHftpfisLNLt0a+tcR
sCO2Y5BZnit2fF0INBOrUwGPntgIB5t1AgCk+q9v+MWoRRiDqvnTTNuCq/RENI5/WpevNxtWqJ52
1E6lcgrbMguKY3QijPxG+yxLlYPx8+hQ8X92Xd/m3Iiac8iwSM9IxlAZlBCxzYvnCBhG5moAwZhG
UebufsYV01i2MYjzub196nM65vbcVGjmIn1XTyJ+aMQciMQOtPw7jY9Xw7mZ1LCxogim8CQuEjyv
xx6mtY/0bcXRpZdkmc8VC+D0bIXT0gYedodpVfwhfJb92fq+wc4eD0RyYdUszzNrTH62EdWPit18
t+0q74S04OrwzJ+nL2EawXOJkVCOgdixxuXGxrbI817mB3VW+G61Utn+a9fc1oO0mxhMm7TqvdD8
/tdaWvELv3k4jcwswKGKZWwzaMNce10Iyxl72McDQ63FqCEWUGSYYyLg9nlasn0Jpy7noPUXwCln
SrMYYMbvh4RH0W4J9qJGafpBiEX0UyXC43ZDK0OXrdhB6ZmrxZcaOz6X/3kRpumI20fMgS2GxmUr
i1kF42g/lO6WhBMS9ju/Y4fogC1zxkpXCkh/PL+T8BSTCFEb5/soQ38Us1kUZHBs98jcYuJMxKUs
+fs+VsyesUH3Ah2gHlCpEqzdKROkkKZDkm9UwrxXjZCpJVFWxpPAnsXBpf8JjByy1yiBpfxawTfn
CKwFChpXMWU1WCDmIi8b0Ve3vql43rU83QQbql7bdvyOVi0/A7f3mLjL4dxbDnR5f498w7eIhRzU
SUYE7DyBH6K7j88QzTBcZMLyCtFNf8UpBHPZuSpHsBmF6Ns6B5rHLUiFXg1xOIFxsaBH1fltqEVu
1dlC0xV1yZMTwIASZYg1Rd69ECMWFJQN4C88NAt5FdIOW1jmeQuGspNHY8kk6xe4oI/7FGDTF7Hx
cGVFnYvJ96cXkEhx3pjy7wN9JNu0PCP7ReNqhWWP5+Ww5zl/mv9P5+V4+gxJj0Lp4nLhjgkkpHH5
KWAQI0eDlnxuartyTq1D5sNGeLtqpefSm/NG/MmZpLzVCGXq8N1/uflECFhtKqIVDLb0n51Az+ci
XTYm27SMMS2auXlGBSjO1VnKrRV6gDiQC6tuX8WmPos0bZPzNLY/bBuyKnLjOHW7W6PgYw0R7eQD
BjV7bWMP8aKXpv2Fz/THzbWemB89bbG9SN5gFmah5Aa4iEFcZirMwh2F9vG767SrCR1Li+jkMED8
8s9sF7WX1AUqueU+wOQYbcikgT2KeafgerjI+dTT2Do6VExg7xlFrwzyh6XR9ZIEUGQmWpGR+wk1
xbf7dwP3nPjX/EwOaw+hp5Ie2JczxGHWUCg8r3lwLh2xzIWo/+r8b7k/PzuGrc+vkxi87HzcDXOm
QCbTPxE4D4Clo/TEq2j2MQrV1Dl3euZF35MnGYIit048vTGAruM2dO7TlkMICudJdEPDn7AYkhok
qR54fG8VSY1zK0PEClkdmJhtumsJwRsFGbsKcV71mRrHLbt9xq0rTAa/57FlCFeLP6c7Mpj3wyfd
xc+yam++K2zVO1zYgitNfKTJl3rnFSdKNyHXmWyqLzdbuB121BfsI8nSvUbxXO4sdOU5cW13FryP
jE6u/aCJ0eOuNkqcoX7qdTK0xxWGwzSzqs7m4p/2Km2zpE9AQ4YjDFzuLDk218d0hSOJMS7gkWbd
pdfz/5QjbiNkcnsRHElwq+uQBb1HgxJkq8seg+0n5GJqhKXPPNkTlwlhTCXkZZKaJs5dCUy1Bdoc
U9gvrWTegbwMzhHsJ6JMSQAbQfUh3TmOptjlfZGPSwJuDdvswJFqqIoItJG5R+mqEjg5w/lCYKi8
VY+UsYTBIm1eoXzoJju2HIiWk27CFUKD/hC+Jk+YLH3NWTv5H1Py0536XKYZkvIJjZ+hxXET5LGC
rzWVCKDZ4BgbEjoRPySndHh4tYIKfggYvUetpBe9OpmJ2kZ7bwJ2UQnH08WrmjKS+eBESigKcdoe
s2O8WkpaGsaAOBXTQmIaVeMAnHVIOGJu3/5Vr+r6iOuzRlcu1O8pdoxwst0YxH7FwjFcvdnMGFet
cOpF3tqBd77bZPaCCbyvVh3ZBfJkaUGVbzTyy7uxzhuo3C/EeFkzbMLR9BuOq36OOb2hobBMpnXB
T6mkvB9dCSVSYDfUI/knor+Hfc5w7WbDm4ZDzdWRcvvKojRDTv68OV3jCWLj4FzNghMcmDLPwdCF
mnFvLUecwtK1e6ACXaCqhzLxp0tsiT9f8ymY5K949XHO1m1jVZywn3JAzifrNr1iIHwG9GChcBS4
p5bQ9HGMLJx9X5YCNB5uLrSrJujmkrlxB08aX7QCM5NUarXGOgoRUnu1WyrobsvvtSRm9Moip5mF
xAsT+skDHBlmiLRb4fQOnXc0+v1P5wQFDu194W4dlZnHHrZ7CAG8NRYxIPcIKuJ+gxZXB3y2NNKw
KXRLiZpummmh66pndsZa/fqyOHDeWw/HrHaBqMr5zIrQNZjSGHx5tEDTbHg2JlJ0vMnA+UGFnieL
DNasAJjnd7LUKppVb6rVjZ/zGjorCLBK2xfCiJD0sfIzm8wcC7fCeDAWU/edb3pYcqCtM2DKDU6v
PmxenD5MjsBSRwU0KvK5y/aQW8O9ep6BwqmjNexypDOCq/5rnAYXZHl0vPQd88xZl/XwMLy4bwuI
hqJv7/uluJ/eLK0vC890KbT0MNOQpnkwVnyE3pWkZ+dsoGSSc1g1DNP/Oca8VbG5hzmO8p8tvDH+
oEh76HRbcAwQv+5eOWDNRDNNoqAcVEyt2WlSw3kKgZx1mFB2eInGvfYHXvIeT6oLJTgI+gZC/Qrx
9/kzg+WyEocC7EfWJFBda0lihc2hVr6N8L2dw9pH/LVm+m+6Yz94Z2Hh7InkaHjx4RljHiYJOcMN
DxcLXZe+LJcwGBsyoK/pkDlLCGYlarvc9P4h097AnYicQhjT/aTGPIE3w+z5Etmr4ERe9CKLJo6l
owyhtj53bgeh8TCW5E7nhQZxusemgmexc8z07z29E6u6U+IxGlt/8TN/L64ALOZC51lSGk5OPvis
c6PdDAG7mbjrSJO/UuhdMWMvDxsJFihltXYZMT/f7Z3+950a1vgD2he8VxeSSACfC4S60bTIY4x9
UUNb5D9Ug2BPID+mek9S2Q4cuMkf15XRnTg+5JWlHDPnGvoNJ9grSoTqBtpWBPQSfJqRzplDG28m
5sTZF2pqypVcV8PDeoSo3mJvnyO02bJPI4ITB8a4gCJGbT/rHXpWRacUV8Mb40V5fFZjxXUGwKVZ
GkmfIRHBSQQh1/DEwVBxhdXg91EVjE2dUZeaknHmvQLzctj0HwUNmugTjNzvGfmqh5w56CHUI/U7
JyeOLZjAs2AHsAWoYoCWpckxWYQ2eTvYDs5roIJSu3Pqu23FHM8231bKit0lUaS9ha/Uu7N6Y1Oo
3Wh9XgggwzNVUcD/McPTCjENZJzASAZEhsuctJXApm1Wt/BE88d3251fX5/CuILyg/X4DmW+oQ7g
sG590jFac9VG7xhTHyVJsw8+Y3wNk31x+cwyFHc/Rrf7s2VmKh1nS3xNY0/tpUO/9TrzfkgYNR9d
xO400U9bHL7xdkdKtv9u3nvtJyGTdxLBrcBxyTf06Gq5GtRrf6KQ75Lrb7SWB56eoTJSUVwNBLls
UaOfhR/dSz/pHikTCOlUZDy5fcxF6tB/Ev81bo2mCz84bbpUMmXBAiFePNR/YxcOcaKjaZyuyCnN
JD4J6XFAzEAbYMkDQxPzIPkESc5KT33c0cdACBLXzO9l9Lz827q9Nqw5l+tQln4dp2mRpytfHWqX
41opo7kTMDlYeok4ZSJ1xZDmAT9IWC8RBinaq0dTGRj9oDjlYtQ59VJcqi3FfJE7yl3ssAD+ti2v
7PAtlkqu1X0pJIq2vFmptUj243S8jG1llPNqG6HVnkq94ijYDUFbeSJ0fmdb3cll9nhudbmkXbmz
TvPxT3IYfusg4yjahmagAVormdwjitn7T1fZxzbUD+dNbkOLJFPJiXReU1Ze9pfmggfTWCboNHaS
TmZ+Nu0QbZaIgm62mGx53iKpIGW7tp4MxUgRuvYnRYAqZ7gXvn0GY5qrb6YNbIJQPJsNBZ2KLrZ3
GQMiWElIUdpwZAtmIpLomt7v+ivPejaZpGPFUaKfMoN5TNiAaITcqe3qCr01KOwki1HVTP6NGywl
HuFPlD8mHr2n+JW+COfASKXmUWHa8aldRF0M35LRzRjG3UILbOnY1rNDkKIgq2Q3/y/f3Iq/JpqA
lvj6QvULfmQ0x+26mvwaKHH6OlyrZUBPhAD7ewaUtENMbA7BiDBcGDnoPvlfQ/jyIYuK5ff31w1F
Sko9lYDm50TUmfUDN9PHqv4yga9wOmum4dLX8NOgNVfKBxOq/L6Ncl2Na5PBYtQ+PwW2AoJxONox
iqQUEQBR0j3aOGl55xxyS5aA7dRDV/ajsXl3wW9KGNp+CP+GdIvakuZQ41D8g5TvvaU+Mg3roGHb
IoXCSmxUxriGA133dexdB/szDIwgdEgtQVRyETjfvG2OXVrbcpzqH6qSGDrdrD7wbmWSkxeA74GN
WFL+nTa9DAx0H/UqXCw4mSdmEcChqf9nYwLILjxpVnTd5meqr/KnYB+0kIR0SUJSDX0T5COYa2OM
K3FuvZukmcAAvOpIc3qKfrMCWV7sYCkGmUxXPtghrVXgn88XMPuU/gBDSL0d00+VI/YqDWQcj3yE
PMfN/rpn+6/gWZBk0+cDV7jE+E3rz5JsWnnUjNgAsN1YTc3XlY3o3n8I6rcZ3XcmoA4eVdDyi0In
Zv8y4ZutjuvmyG3DIvowkjVB4OrZwpnAfu6lF7exnuBVPyQHmC02xU6cF1tfhIq7+ReC2n6eJmDO
2cVH5FwRo8Ddsq7BaeH+jfwVj6S4jivhXwMl5eU0KF22tziefL82ZytTOYvkuOnlCYxlIkE1WrpL
dLZ3fxCcgJZhSFIzl4I1n2boVIY+9qR8I3aEDz/heMmmkJu8nSQz961Yz9Hpe3u5+a61lp/kE9r9
t/3e8IXUB7ccY7V5+aLtDWtBXv1MNtRrEoXQG30CuL6oo988fYeEomJhMcydLAV57SHvbgWnlxIc
IWa1hSuBktyLmxa1fNJV8ARY8ZVXBkhkORU8XQ2uv446y6hp/CW0Kce7aBt5nJAU7o7iuWG7Yf6s
qxvrqsXydkJveMu3HU5xfW/fyTEhtKS2jipXNAWTuP3Xs7+JoIFIc767o/5K8EOXGZpi+NgPVzu0
wCLo1T0lWJf9W2xBWorwnj5a4IHrsL5tCir1m1enItUi+sxV44DhmRmmSD1rsxGVqD90lstv1H4y
m2RtwpQ7BxocVy0vOOuoE8vR0okpQifBEb7VSBHq5Dr6LqsqwbYxGf7623DtZH2mp3XQRgxTZnKW
08WA0zDW8v1pnv291+wR1CjdMhCcLpDa5n515ZX0bak9ylSWaZ53ehDxI67cudHQ994n9m7frVLE
wuQlgCK80D8nk0ak3Btc0vhet3wFKCrvsVTJ9b9qHB9lJIflh8geotvjQEZNfT/x+0SLH+pmFDKZ
v0gqhKxVG0Rfw/ahnodlqTdfZLUhvqD9VmXRvI8DGKRDXlBHentpgP1q9WznV8TGcKMY42qSDhAx
6XGiXsZj7SOMM6YozMUSMqKrX2lWnUIdIAWICKOeGHdgGP1qTIVAJuyPncMkvtx1trlBlJYTXF1i
4wrv1gJgS/SzQbr/1OCMDA5KWeATjqBRJiJBX9YO0tSDuWwlw8hcgJg+evwwgtpWaBTk9TyY1ciR
sScP9AP3h6E27fg3RpziE/x08EL37Npu8JeSR3W2F911Fp2Zm+yU4I860jorhd9XjrzsU03+fhOU
RUV+E3LIE3zKaT3VLv0mo2x4t1mGp22QMd59eyHmebn94a6cnH2tVHSYwCSBAT0NX3iOseNBQGwO
sD4/tV3O9PkfxsQneUnfU879uTsb++Kcmi25L+OdtvJynJm7IXWLlbAuM+G8LF8kG/HUHbpt+9VD
ity36Ipzws1SJi5aOjMgGQ3MFxPjz8kDCu0OwJQr7j6wIUhPz0eufBkUjhk/f1FiiZGXY/lTHOEr
4yURst8pMVWmrUl1iCwThVOlEiOhomlej8VoODlliFwd4mUmMo5/qe6cHS5g1QzOgK/B4HFEEqIS
KBNrQ9wRlK6EWVkFXYQTZRK+8y9Ed9RGkDSsFYQ5Hjoy7kNZU2M0vYo+oHBipm510++NYSonuofq
AoDrI2dJpQaGqx8ZeXh8frgO01YNH58Jh6waP7OiMmyC3o1a+7yv1bOuH4vcRqszPNnzoMbmGMN5
4aKEECulFoPOxbYCNF1mVweEX/f040wVHqXqmVvrWwqs1ruCKe2cI++pHZaNx9JUoMDofNms7kFc
svndhdyUmSyqHQ58nHFEMgt2nPX5OyHY8RVS/snxwHBK1G6jvo43Ol2p9EOvQaVkb7E4+j4YPc7Q
vAPhv5D274XgeXkbDby5Ag1ygg1AApbhwmuiy3JHAPxNKxEoRaANYvwZ7Y0BINBk0wqct6aht/4H
PoWv2Dbfmuf4kiEQeHjTOCZgaRXsXRnFUJRVPKkpBvR9CHcEAY2SrxpOamZhDMXV8lJgyUVUGOmy
IJKho7IDsV5Uciz6GMjaEo76VT556ZdDrWomCjq7a7c8sWIH4QKCJhISZ0yX8FLP/duooEAH3XME
NaJSdQQdK4OQsBb4CCMPWsiWZY1WHyX5mIbuLsfJ350iSNtbZeE5YKRSSpdrXkmPTVweAbbS00HG
DulliC38KFhkRH9xj1ZNkGxZHZ+Ku8EJQWLYJbCG4lPRD2uivZLkBDIH69sCzD42FBWwfDIZH97p
7pjGd6RGJ8dr9Xl2+wHuTywFoJ2ZNRQ2gyMJ8NurJ4aE4Bw46UHkPYzhXuk7f/v/BXMD+DQT53p4
/uCUOHSZgOd7DNaNQV+3M/f6TZSlAZHIltWYRtUP15Pl8ckXbFYY5HYyJjeTsnxTfPSg784OsHwj
hsIQCzNSAZGRi6oAnO7lLgXLn8lcqHI8c0GxvpU1P0ruNELZtkABauYmrgbojDIlCo3RA3OzHBLE
Ccp81WIT6uXxzBFKRTgDTy8MQqBZlpVxVhOeYy98Syd6YPo1Os3/E6T5DCNJXdefP/ymS/pqRgxr
D1uydPgqK4YngdlvGeNgJ4sc1ixpTfQsfsXREeZWpGF4dKk9tDO7/7DCUnyDYmr/8IhUjp/nKV8S
S2LNb/btAH73J7gEgTbViuvC53irNDiOA1yAQBFUs4QOyFfBgWDcJVAewYMuhnfCXelPyOZ/bPAv
pi4GsjCPXqxmOVgS4OIs1rwIFIN7G6mO5IcNpyfdQOqXGD2e3jdX9SvlDLIsiYtxwU5y67L4Cevz
qAoOktcX6P6tNRrSz9l/FTp0BUy4EUwbRI4ih6dQga0/NepZvUUg6/lBxRjmQaj3cYM+DvZKuXsH
x7fTmHTm6zADjo4kQC9CQAMX/2FlBKGSM8hrbunpNPw74jRi9jT+WDVF8fq/01AAGAUvsMBbzDwn
CrPybwxNa0pn40lN65jeqBs0ZBemMMerts9/Min3lu92IX2QDRVDwtd6kcMs7Av00Edc/KqaKMf5
hZvZsr04hGW0B4lW/TXStQlAUKHxj6LSqHU0EjLgbTbYgHQMIoRIBpxSFASBHggt9LaZ9R/gMmP4
kJOQzuPCLj2K8gU5rbWMTAYM/5VXkb35Eb02lEnBKYqGxAhn3AWTCJGAHDo4Ql0wkYUz2X/dsz03
404BjTt3N7EvJ5Li3nYxMKpbNhvVqxdnPhfY7k1c7EdxD6+RTrwbS6c9a+dYNbEusO1MvNsAf6yt
mIQV+E6xB250vaX+Jtawsddx1JZGsqTrGer/oFBQLmud6EkepzHQG3AX/wGL4HqG13THQZTduj3u
7YE5li22gcp2wy2r4gDLfJvo3TA9L1Wp/ePuQgYc4bD3pn7Zter8SeXG44mXsd0FDVsbWtObCtDR
9fm2ieGfdmz1+/b3Q42Y3ZT5MBYZUS+w3KMivSFcFaSQ+/ISgHU7GtRHjw/UBE1AdgljEmZ4r74/
0TXSr0aOzXOpG5BNRQtxFhDgxZZnNgA6AzzZgcsoITuvnBuix4RgVVZUUVl+iwnbHUYhd5hPprzD
lzUbH9kn7Lw8h6D3dngLDnlpYnlZc12nO6ZzReN956MNN9oGINDPZ4e274Xa+ofLL94U6XdhOMDY
RHwAB2/PwYcTR6Fpw8J5RrJcCoVpngrukuCXk+LKPXJuYbyDBWC4tyU04xv2rjiW8tptWiFbXHW6
DiVCt77rz360RhhO3GYieElBRJGSniPEWZ7/9jZWwMQTF1t3TK8DwrulviiNjPgFEEuycfEfO1DJ
9EB3pxaoIc23tYVcDIT8As4xrBkjdKdIRz0N4DPCmsb6UqeG+4Agmy76Ds3Dr2iT3MF/+QZ5bjfD
+uhbLDURavThrVkcQBpXlSscoZfVIoCePb1uaOBrshEY2TT6pLbqUJg2XolAA2li3ixyiWBMWhrf
lkcWjKmuL+MF5qYVRUUlszdwI+Crv1uD9yMHRZy7QC+UsLb9r3/x4WksVPLJUFx++4hs5LUYM8Ez
lvxb3jy/F9d8CWW6UOn2FFN+E8tb5pLTbqPePaPmZWxsU8fSf9tqHcXIYUWjUfftE/BPbMhuQtPt
rxNq8PrHeFMNrzNGlHGh2S2VJuPCcsPCngz2YcZnh0aq0EDnxlShCfIq1sXch2snAplZQn3KVzk7
5m2nGp6EjWsA9pTSM0etd4wDgsr5BcUKXfBKCPYFPKL9Jkr4b2puiKu57H69xIO3hjDnfT8/umod
KwXKiSayTVnBhjzMATdGpP06G7u+zIeU2QAbDMp4SIUU14TWbHFQcu3F74subo8rVGyXduQvFgh9
wjtwCCcz9K9mZGVqTnH5HBoFrKPt+sk7JMH+t+JkR7pgyQm0kUyHLj1xuO4iMMEj5xqpHV2kyJqA
R6OLlZkLaU+yMfHmwJhfXqcnIcfPNHA9DOyj5XJMbwhuFIHq2tAaKWaooQt0yE65/MritG6mK5/A
DngiASZq5cBV/UYgRx4NBrTLYWakrQiBckxfOfHn0UEUt/OA2Nairgo75IIpePPzkvNb8+VYyvwo
hxFP0tXgF85/XbwfohhovhWUYWUWDMEAovFwbi8hIE2/wSZkddhVlsICz+ORmbQuKmSUf7eodKpu
GYMtziX0EdrSnv7INQWEvAxXQ6mL+cKihElO3EYrYfSbbyq1W3rjOJ6hsWBaMDaRk33xCAf5dngw
/GgW6W5fjD2opsOCrZ7RjmIV7DHofYa89VZuP0CQAAN1jhBne/Wq1y4/9evFWR0QbW4OnFjU3MYN
spQ4rFMteKMJVjZ+tBwcayniWTKjgpMuuUxUluO3OJBpixdvTgN3kmlVNcZx05SzAN1oMEgEeyQz
F8PifqkPUsOSQGuByT/A8UHV9Sb/VpCXxjBL4aH7SEqR10rVojVLRR0AHd99VRmLHsc3b/e/8Z/J
STvXfJHqnWClcoCm2+a+zFz0UOf1pKcf+PavGtCIuH93mMKS+mWwvfy40TmaAa4P8SwShUfE0O2p
RKRy4NJEUF7HFq9tfJ4o9FXrYg0+p7F+qI1CahXMzR+W9+EdNvsewUCNjPE6lFjPYkgQ6SXiimgo
iVX/ADIE8eILWINlqDCviSjO6MDt0KQktiSvAkkqfXp2MzBnLSrPdurnxdK3JamCpxBQSPkKQqJ+
IrX7RVj7QOm32sx7LqtAGqstLUmnG9QEx8Oi50uie1MIC1PVzr+XKIM/GK4f6KB11uBFWdf1fg2S
2gnjDaIXGwksept8SRIhZCK83u3G+ELQI4tmLF2+jmxsVinPgTLL7/e3i6b06A+TC0ttY4KnF5/k
S8SmqZr5T9ShIDN5FgJubdZhCFTLjk2vWg/xAkpFDCiuFmWCiwuzPnVT9ClvrjjneikGo5jVu/vf
c1QI1+v8xv1X/6L1bE9i071TpJLoUCRrWaACzMvSXZRDVy/A0F5SYIj7QlRLskcCuuj+lPCwhZX/
lMvM2YrmUl5r5Yqcpc18Sj9Rs5e9hz6GmAW3g8omLea1ddTpC5mWk7fU5HTxIK07mPD0P1SKyFPN
mtEXk8upcSwovwpqB1hjXLnMqrCC4eecMkwCNJlyh+Gc2xdwtf2EmX7hr0iw59mm5rhI+fHgMzPg
pE5512GKMxhVqhegH87CUXAcFtttQuiTXkGhcC2iluPTNuvcQ4P/IxxDRXVgqZQcrU1DkLsIe/v3
24id2msnj2YDenAzrcSrR4+3yRs3o5Fq6/nSSMKlBF8DCLS7fXgh9trwEBgD9fa+bwmoLRfKKrKE
dug7IqJnZ+WWQXdI0yxGlMciivG6j4ZD+1Qn2JiNrwvhl/Lhvp4z9FqU05BNg1zWHq5Jmgbu2shl
WGojvz1FyuPRd0ae6FNNRWvEanEl983vbwjIkvntxBAKxQSLXc+A/tKb6J93qjdxu1jXo2Wf9df+
UipLPgv8YLYIY8jmC3+aiAofWmDUSn2gU90rW+Uf9y+SCWXfmxzzGILX0c15ETO58vaNfVUeITOw
3VKCTJLgoHwZCBDnqifpqyN3pCpRrgUzYPLWAhLa9//VsNVVA2aMWiAUPu02lj8M+ABYsYJ7DXaO
w2H+hbRejTkOn1J6J1kiZP2acez7K/d98qh6nv78sf3gUVEVwe/oogc+679hU/kYIdvDAHoWEDmG
ko8RuM5+xPZLOjInVcvW1cp92Rp4O/fS1qTtqBMw0PBi8NMw9ZPQDN9zrHAubUBCxOzgUTc1CKCv
frTcJVSrmRrx6SvJG6BNzOwRXwpV9fbhJnehTfSktiJ7EQ0D43e7hKg4jxTirQKM0ebkY/JnP+AH
KQE77oLVOaexdy3ycBPkfGBl1cVC6oQ/9TJvdgPuiaGkudLAjL5NZe6LwxZsIqbom9/PcKTHj4qK
tvoHc3NojXM2+a0O69bsN3iML39ftRDNlySTwW+7+jL3WU/Qyb6NG6oBWtrKps/5eGqweNtczmyE
j/0QTu9HLAvk96JADT0QfhBjUL/Sm1znY0POCwx5izqntkD7zkBCKnYbkD1LQ3wNs6u6rvceoHuR
I0f9bVagq4ykfKS2pbw2OsM0nETWwxvUH3P1qOHH7PqGVDc3z5yX7t8Ste7cPzH8CizSBxsCNpju
7PivoqH7gG2TBl+Qi+RBWN38nNPmRWzCTl9IitzqzRFCtUfh2OgRjWfPh3is4f9J7YTIJ4rQiC31
v0sNQwK762dTUv+rJAgm826+Kdw9xzOJMiz2dT13S7RmL4YY4H/EjzCuMwng4HLbOHMm5TF7hI5u
oNyAZPSJYKXZ8TwDrr3gHU+nnxLmGwFELfdlDHCCjmmwbX9DGMO6TWxODXLUwTATz+F3G0UzPJBB
TRkDvXEhLs5+wEhLvYfWbAzV/o/2kamZwzCS5GpRopdXZM6E7VqIGpFbk9bx9XtQiG4fLlr95S9B
QjsMhWGXJj3BpSLYAtBmLw6mLJB3QEmxunUpqRYsEWsm4XmHCALNa9kDaC42HgXmVVxk6DCWjUQU
R972KIjQslRlZo+sQs/Bkf736asKVE+OM+2BuSGrgI06YYmgcQw1DLr1tBp6lDP03ACSHL7IByB8
0ag+Xe/IXYY7XjAOmOzblSi6jdOxOmfkWGYJK2uknTrNtOrHmSr8Xp9DIBwE46RFwOa9q8tIoXVG
eBPuCpRKXussyn9lhymwA54JwpvuNWLN2XBxV+sQ1K6TvSjHgSXnJ8TQVTSmETQrPlACM6Z9BYYT
Lood3tEdlMwQM1oHX0DZwT5rO9phS39f6vFkkWzZiotUadCAvvvIL+vzblT7JVyUG7Z/o3mb6T9h
FSNPevlKda6rRHWau81gXmkCwUrXLng/5L303VVnDn4Tud1ue8vaEIe8BR72x6DIiZWmHLvWwzRF
v4WsVdobofaf4AltPPx6YebJ7C7m2hWiS3PE4euVMY+0OoVVeMMFJe85hWJ6g5YtpAkHSsL7K0eJ
j5tj9VAdcdvcD+FXjej5RQJbWLo0x2Pkoj3nTAEXHafJuCTjmRs8fTPmzBcOn6QjorxjtcNT2mfk
ewz2MxlJP1JsS3dmxcHoKr+Ktm6JE+rvoRd1pG5V8shBwURwGnwgYJLjZB48qDjLPRqQRoWAXJOa
0FTQ2HaXLAdJBDwYrO/C42Sk1kdKLHDA6Uui6CAaqQ3X4dTRbwCQIQbsgsy5LV7QPMX3fRHbnhZD
pidi+ovYG1m4H/sU7PFkv0labUVbRpmpRA7g26fhYmxyxaeNKeS/2A4oxpTsAEMvINK+sh4u5Pdc
LIVv6k67jYFl5SFb8CtyfaunkyiWnePI+05xkK5tVoA5gMLOsZZVavUuT28yWW1ZUMhvS5poN9wJ
78vDYx1WET5sgioW0ItYvwipag2vpew+OATgrL+oisjccjl4W4t8fX+EIQKm8i565ss4/zsnMCTw
LCCXjBgAToqQuSkdRSy3cOaF0iWs26i9HP65IA/XOpF0eIlxYvnx+L8FYteYttUJx6NEVxmHfDuK
WY07SbFU4clG2jGCsAOQyJeGpPKIpY2BgN+NMXFCYow8T8b0YiIPmLPVHqrdvockgT1WNa7+5etV
GcYOkCv7Hk7mE7Vl7wir/yDk94qsQXWh6DutJVcKdliRjWSqMR0vKg+S0nWmeGAeFrQRvF1qOLgr
dWzF/nABAZmL/6B0QHClWAnfyxryYKY3lK1iVJ3mAQpXcQCz3crQPhgQ82KLNBoamdzzrY56MZxV
Zv5DgKlBvuxxX2+59ocH+GpKIPw/Yr8ijW22NKocCyogiNOlng+mDLdkxq8ggdEwX0YZ0huywmRW
XMLj8ebptXU33/6e/rptVEBxx2EDizct7JLz37F3+/QcMgmeS32CopZEvrBIGucmrWWWanZc3VGX
2MilQMxwA0CcZgK1OS7LSdlLS28jPMN8sPi80VfMAyqzX9ZRjm9nbzV9wRAc3mNeLdUfeAoP71Ht
OUxLbbLnXDutEFl49Sh62fwaDbs+gIYjtqB6EgNTmu3gpQnGQVPkE+fToPvKn7clRn2AxhAwW28S
ARXB+/A71tugD+dde7wLfyDvYlY5n20euHpp0+DupWWFlrLlBuOL5r0OBiR4aoxhLOHYv1VO9Em8
Jqt/82nWyFwJPn+N1bIYTc9KbGuCPGHz23DrZ7wfzLOJmyLUUIbjdzn7sYyrNXm+y3XGIluzuhoI
2jymfGr3vnTYAyFU0rlOGCS5fv3CiDkwWTxrSSiy9oivSAM7vcPwW1qzZwJc6ytbg8ByemOB8aLF
PuayjA717bT8G7jGMy/PNqnstwnY3TtKsbZYYltuGowhdlj1UiY8z4Gd+5pwmeFk3IrQP7yFIYmB
CgfwoxIDrVqYBEFmMqHk7go8d1TqqYxc2HanL6ktGHmVxhdIfrtzbi8kzwnaFgywwvAnwWQIPpvt
zrZUw03F0ZhXBlCnitK++sFw6z5EFVkmCnYCnge1tH5X8PCjglaNl4j65y+oJaK7cfgA2hs7mQaA
mzIkbZgVSmgbSxmo+OrI2uzeAZs1QmneiMbrtP7LUmLwg9UIh5jNjK6Dzg9R8VfhquCAHD7XF7u0
uENTwuJPLpICOmRfY5RZOBNq1Av0KvRRQBHvvqq02wByPUg6WK1Tr3qG1NEJNqEVWCV5gvm76H0E
3WfrX6uAV9msHGnZpE/UoxihdcUmXsyXq/lVN0XFu4u9jWNlV8xn2BlwaRKxMORCBLp6DeH5YR0B
xUA7r+GIU4r0aKkmFsIA9G/AYS+KE1muh81+llRLh9pyT7RPsvhipQPnhhtojCVtq45RsgiD5Azt
BmbfUFOQp5dvw71YMtNIDg1oVE1uGMoHDSVwoiErRR6lIMRg3+a1CLV6cP6ZWD/xsWSeHKOynx4S
kfyqDQkqtCwlB+gQC8U9Sb6+Ig334xUBGC+TUwNXHhAUsUWjy7c97NC6NhJb4jHY1OFeIMGnaL7S
7GIba0gDrHh18k0ShA7/O4iegBSSbkdZlAIkqzwaOpHWomT/Oi+7Q0cMpC5owdx0h7hMcxv8t+GC
Isu0FUi51McJYhFm+4CJhXlbyW/x9sXTvWP1GGODZBIJUs5wLuI3tixYo4DvL7eojLCVC2+lKaVF
+xiuO3MTF7jRRWgDJUMrSYAH+3dqfVw4xlvybxm+EX3s6qRfzgy+RKk4NjM8wxblER1TPu/m9pbT
s+orwwfbzbiKPz4AQtar76SvYv804unhVJGj2kDiFUvKmAiWzVOR2FO0ppSbAsrmkqBQqdyaIZmP
Z3F4AeLoZfqZO3+WsQzR5BxHwscSf/OSpDmtjo+S24wxX3/SuISLU+lf8ECrjU2/Q4az0p4aHRht
Xy3G9A3U3xWBXGAJll4N/esA04WlxbvWBhqDbSpq6PdW60Zi4TRe+ZhsOtXTXDoLGgKcifV7kz6o
36OoGp2NahmOhnaD4mjQf+BCc4a0c51HhICBbz6MK4Lt2F8kSv7h+Rz8k8zNyIJgjhaMTlDFk5My
eq3ONZsuRovE8d4PiYDWdNk8bdt8W9bHS91/SrosxGvGZ0XpAWMtjJ3FltenuWNW6OG/91slihR5
BPNVr9sLXzA7PV5y+Ac8Mp/ABpAqb9QHwo278NCbUFR24RXBXkSd71Zhcr+FMqQDsuT2ccQfVvGu
hVXnwU8EeKLtldS3AO3QYKtkFqdG23BsmD1oEUVJQPa+NjoAxCpbdVSNIzD+x2Sr+2Ccf5QKcHdq
GhtVo1ZBGqAa3rS/vv2fHd5idIReOHaIep8PkI6rPynhD4ZcnOt0mxyFaOlJ5QqNy2hnAPXzIn4W
KdWcg0QN1Et6PSD/EXQsJpK/Ik2JHwAeigzOvSuW2VJukXEWFvZTn0DdFChWvQ1wSorrqmnWLJG0
WfNCewDu5y2I5ZyoG9sBALc34QJxaOtMfisEO6vmYKFW+3kJFJ5t9c2Htp1ZrAz2Tn/4dtiZYg5N
PO1xLCeSGBdVLxJaaXFQPMm38xMQ4gSsB2EqiNFRoqllDytWHNCgiptJF+uyf20MMlTFJdXJDWAp
gEeMtggfCnQrQLtGcFhvqr8keeDx/H7oGG2LpScMIvMmzRH/39dijXAbOlS4HG3l8xgQwvAYsex4
R4jrRd6UVLVB48qgtW/YimhPoVIUvMDcCjjwNM4yQSRVr4We98tneLPNdw/OQvC69ikH3eKbV/4V
Zi94BH49tLgBtEYdtQw8cIT1qWXcIBUqtfYfAAT7ldBPYPzuqSCPgus6hd13SQtpZE3sdcGREtil
1aK4R+CO5OVXBgMYD2Mvv/fJDh4xDLcgoU217c0j+/KNXQbFRu0WHejes4fIL/qV8z3bk/G3DuKz
G64+yXLkxmUCJ33tZiQc3ZrPhQAQaHB6t0/lLB8wHAxWEg0+YIMpk0IwdI404kVooj7X9Z8b7Gcl
2WMSDpjkzq5up0JnfEXUyvvDrPqyTGf81DGfnWMK/Pb/El73mx1hyMjHtUt55Frqo2ANQlCIj04X
GchqrcRMucMzNTHrggQv8T6Op6taMKJPRASMWTxCn00Mux6IfkblQ/s1nJR5BVLi0h5J/0k3U4Vy
3rzRffHVXeWw5KO11B/lNh3jnHXTtEBq+4iBqiRq4f5eUMqGG1ifOrx2+s7wHisBxrpvHSYNKIyN
xRaN1tk8tfWWSIn+egolFioxFZyR2S6DX4c93wCKulZX3A9jbfki5HNWR1UUpWvfczahZ7aa+ahQ
VSfsnLhR4Vb3dNQIOicQ/YARPQnCh5R8SE4O+iHq9lDjzCRJem4u0jerVyDHiwQ3juZy1lmgEL9w
gVyT71iOZycsILUhh3wjtIyAsnasy4JeV419iLRkSiuPo5VoSwVO/a1Il8RN/opm8ayxwNE9kkSN
jU1UJNSb/cl7b3neRPvrZskgEXuakZ4nELPpq76vTJerYCXUFJaLb6gnJginszJ4atbZqQVr96z7
eYGqOqlno4wclPJKWQYvgpMAvrvtWUAq4TBXGX+wkn6+PtcnXSRfFlBwEyvjiSjHaS4IZWkByCET
hVTIMTB+ZR0hEG8ztDAUATvbJWGi5bwJS9owNRi/huNScyHyfu4TSl0vDvrxxOiXW0mguijhxA42
dz2MnrYn1p8e/KFylkUTnFkIXeBM8v+mrRz/Eo+y9t5rMNY6mwt7rFG4VTfL3WwG6mEGSE2Yvq76
dMx4/rSsaEaQH5eirxVpRO7/zK92QL9i6R2h8AGPHjf1WfRZmMueELSU2DjlrlJHZmrTvR6RcWya
gxTIRwq6CnxOGLUgNUohwiT+YRUPOldowhDUx+LTwN39kkk9KVa+rWnlInETsvdu5i6Kb3adSD5+
gvc2JW5gREZyZFlTBGo6cwyTcPJgmQRvgx2MKn691UZjbNzl19ucYSvx1nEZQxC/iSLshmlDD1Kd
c6tPTSoh6ifO1hKRrWGBafW2+Sj4+Rl3L04Bpo8g3Pestz5OTRrUOspl9PpWBjLjXpRQAy0QfKac
Boi/5R3RzUeFdWM+9vHNnMWHx/+cBqla4TSqU32htDDKJ8/lIoty9olWh6SpiACgx1QNGVaRj8n7
GbpWE6N0NkH2WAObCA4aCf7UAwBQlBEj0hMNL9Wi25t1lFqyoWMHxgPBYUamy65Jxe5P4lOsHH5+
k9GYV8+j3GdCLDI21lYdck3+TzPSoqTL4moapY2QyoytM3W3gO7WoJviRLYxHQayMr099IeZH48N
3z4olaB3X5GzWk06BG5bNwqkur5trQrraT5Hk2MCbSkRG2eBs2WJoMhp3F8L6rviDQd8uRBh/9wR
9ufq6cHgCAV/WqR6sJSeNd1rmiq5tb9BidwTBu+AdPsVDDwhurbcSA6pS+KuT0wmXbWFBJTaXOZL
Qy72NK5ISGwa9Nos/KVRr+k68Uk320uWo6Wp5/JC9aZOBoa+k1H2DBg+OEUaLZ44psjThm+c6Flx
mzYh693opju/Ttd98AA0ALun5dS1c+VKqfgy0iBgYBy7dJzNnK6+eWsiLXRupdMX0SmpcxJ2NvQN
BDdTZ3XqD4KY1b1I8DulzqiqAc4UMXgwW6Dn5OxhTzwPfZWU5KJGnQyG/cxPqFr0LjwxEg+9Nius
tnEYt+LlQu5cGNrq+5uBwktD+MgqBBjVQPjXPuOFY5jaNOJMfoFgrRHcJiFCDHriwTAO4tE97vsb
NFvUbbrKBg+MnOFHKh/s/HdgYdNtKf4YgG+ouoEgcNJL4biA1g93nXGPNlK1uOr/F4DvzxyeYJs3
HmiCM2kLWoGPyUNKNFz13kA7pvMczKutIQj8HfAdY4Mfng1CfzhuN5Vr1Ec2QSH6QDxsZKIapSTd
4KDKyTRC2c+nqqrAK5pfTBXLqkqm8nmMBg8wXJo2HUT9AQfmXSCp/5RvAHUQ58NHeExFeSwsWU18
WIQ+Pwsf1sHpc6S6P86dBnpQuqriJRt4Xqj4ItOezi9oO+vLGKCKUaBRuLCEdbuuTJmfAVT+v6EU
6lhmKgDukC59VgcX2IaIn7bXrPUekWL0gxE1rWVG9G+fELZV60jSk3kaIfc+3ZDVRMoj1UMT49j2
wL17IzYGeuvuj0u3+AshG82ARu+qnQXFX5p3NVChvMK4E2s6De7ncjLHfCEtoNL8onDt58c0EAEB
udlqcHLfPBDaDccGCNF8mY/xLxbY/HPYblc9TBoDgF7cSKqy/dLDJnn90cLemDh2xsoAH52N3V1L
0AubSJ1kZXlsfxHU/fEtJuOptXT+4a7qQAlwFgcKgoEzVszhakVwORxn0FEGYksY8T8EkHoqGwp2
j6ZfA5M1sYQpcIzLU9Raguri8lxVm9I3yOv5nhel2BrquPVwl4PDmXwy9V15UhMNcd2W2cRsy9Yo
lG6EEClEI/tfOiKmFjvjHiqVbgGoo3jvf5M6XDdLO9pYhZ7wCO1Oqs9uD56YEWjiQVZ8WZQ2szB5
M5g9sstgwaIFEn8sO+jiU8jaTfxMNhHMZ5byBSAmjzXWjNoZZ8SUlEJkj6Mk2ZDMLFFfV0Hdl6t3
knyKSo1MsbMqSP2gA/6BnARLFRFjtKHx4Xx/SJvLZzrpISVfzxM5SGzUGlRNXUbJOoMunxvSV8pG
C3HSkv2TNVwWRT6oEDthYn6rtGCcD01VGGoe3377uNaaVZ2MRjIepz53SJIsYjw7Ob4Hdejss1jE
IwKcmg/RsyXTIp/OHJhlPOyMz9A6Eiipc8WkcWlKJKSXhf64fe9I4c0EnPUfR8hPljcnzQ4jgOEG
ogOyssPk8tPrjRWwdKT4v7eKllBNhO8JQRKp70P8plSE0v2lIGQEq0aN5z3xFZtSYxrXiisNdL/N
yS6/TBx1U+MSom7rUzVoJwOMXPYlNKmFNmlepRPby9ygSjmVU3L5uAF2HMqHUya33frGXmIqRK3B
gjlPW+/xiZ/IAtfb6RLReyCwhZ3MFZkazic32VqbnW0cIZEYC5pzEptYI1NHoSv80kQ/0ENp/8SX
IObUJAcQ93zAbpQfUgf4wdar5gpFA9g0090mj3yhKj//oMaMpJN3uQoNReW7YP9ZVmxa7umAJOWe
UkoDil3HA6jtmCasyH1VXyljj7I5YuPlsLopm8+QO26dwm09IJI24ZwqRjPFoycsL2LNhwHx/z7i
MWTaAo63IREHpnXy8wPy2zWy1K4uvWIOV3isD5ZaPw8aIbZmYSPQalQgRgSxZzO0cjv6EzTbokGT
h8vFYKLJg5LJLgEakcH9k0S61V7d9DYjsuicz/f77ERrsWPf4zI7a4ksroVOxRIbEXrn4x9tie5y
k6J9TPMybNB2FCpdWas9YMBa1yrn+1v71MLGnb0PvdJwIwrqTDpuRhsSmX98F8/eSC6ho3jFOX5C
rl48mnSYDGoLNPd822sV2XMTxOLfmetOFqHni10oI6urn2H+VooTywgU4IvIRNw1EsiJUaxH7J/E
Gtddfmrfn7j1pXMc5f8I0wLfy+cTe+k2bRhD1HD/HJ6ri4kgjS8HLNPUA5ud8oy/F/VjkoLyOCkl
VvrqqiHMl2etEXjx034jHyVISF3KLhIoDPNB6JT4SBANHM9jxAVfxfelySy/T3QnHNlKfzFPYxI1
xIBwfQKijS4Auc5oQ97Kk7IXierJ8UrCoS813aTwwOzuhWArYyoNQjoT9J7bpZBLRHbzQbQg7GIf
qzJUSDZpwlVXwsySy/74wN34bqHLFiAjQUsXQ7CD9dCI0gZMGZ5TNTXXHBdsPOMZBiyqSVfwinN9
0s+kxvRM9vHYp836xAj36mMoyiLcPIkt1hAFr91NFjeXxsrrTwHbVHwEcVsO2FUM91anOzfDdEay
Kq3DqwFUWt2A4TJ2HBeMHdYvqzuc7RgyccOE55i3FtZf5CMMZBb+v643sw36ZICglQ+RUZ7/msTc
LaFY8wep7bgesWgK0cgn+g07Z0SwQcaAB8Ds7MqR1Z4Ij5GRsk5Phk4W2l3jM7My+sEW1Gks0s1x
dEWFi/t7BuLczJ614GAaRrX+l6jGtsT2b1K1EiZiGL2wtoqtp959pkyTH2wOKjA+SUFzO+Oj/Kr9
BEVbnWDO2AdyHM0Idl0ZQzBZX7D2tgmg5UVRwvD1AfwfONXT8rWXV0331+vDumj4KI3sQmxOchva
85QUjgGYO6NM7CERSAcGbOLt4462uOtEJ1lB3ktt35bB7ZdzIaSnqfWeY1Liy9VPFwb0YMpnhLv+
SKRChAeuL65Jp+sKFCEj3GKWOPn6FIg93Tc8qscwwkWV0O0sva0GNiNV999oM/rRgm2C/1D9ANzc
YdCzq7WubLNRiBr7nL5b08HtbsCucZ8kg+SCdMuvX2d9n/EJg54f6KZ3AsNSel3/Coppey7x29cC
ca0xEXTV8sa7Hipq5Bi2UXmVvbL+K2pWpPsh8umD+HQYQSRZ24jRAl7Ias0aORubWObRgj/wP+Qi
hnS3t3K9igMit4e2m/hSs4BeL4HXzn+4X0T0kCrDyeQZFU7Oj2UszSHhOd8j/VMceRYpffdAXjyu
HXmeEWXxY5Ny3lZX/z2lRPcIAk8fH0TyMD9iiNwNn11C8q2zsLrj5p2BZRyeJMseBbXM0NPkzC2L
Tq6Wl9rt+UcC5/ynKK8oaJAxPulDti25oInV0zhUsb9mhZKIcQQEymBQlrjSTGkm8gBcAoiaJl7B
wnXRDV2EBrROeGVDCjtpXAFQZjT1BRxTCxhr1IVTEe+yYkjJIXe82IdsXpsxuOhpiBD8/L2og0Gw
tW/Q+njj8KSttkBMb7T8pipPSkeHpS1EM29X+llfHKTic2n+KsSpcru90BpLyXbIRLEq0L8PwQhG
uCBGbixhkqe5KCHzJ6JGWs/B8mphx6SROtGxQmOQAhNl+qIBSsAs7cKpRzGpHrUtWIQ1V3mzd1Lf
CrlXaYxUuMDsXJQDtUwbGIZVoqYk1KFEvaB8E9y4Dhw/KddDJgNzOpAKS/LXS2LKcJp39EWQLUb9
lw7l9jGfqoMHzXEO6mtZcGZzHk/zGqG7m2WhyO4ZtM3tCegiTXRlfUgllXK75M9vV1g02aqak2XI
qaM9sMHdmUq3IPLLazdcK9DSrWcHxBM6P29BqswTLZQMcR7ZPnoZOpXZqXzTs6W5dp+Rdd1ix8zM
Pzr10kDbQfOEYCj3jtpHK2Tr86GvqulaoZ52032qAmmQxUc5Y5QYdjr++Ku20zHmCUj765i3OOQR
UOszLx5neLlsnVcQ2E6q/7hHNqnL05L5+E/1L59iFC9OE5aVqu6UjswIIEF0LVajwESHI7Eo2+kY
oI7Dy9y5Zl0Jo2FB0+i7zxnBqUIIwK2t+lf6isSN5uvbukN+GfGnU/H8FHwSkcoXu5rA8Zwlswtd
sYOhMxWWJ5gOCNVcL1PfFiFKRn88mXVLW5Sr0XR+ahM9t+1l/hvFqKkRA539CHLlMtGbPj9N8CL6
AXcFcQmfNvZbwtOW87FgWRrBbEOWcseQ5q1lqEerVwgUUvkX1YkpQNvrjNf17P9mx45ap18jt4WN
opSzlkVyKcwNGCtowgnt0uv0LCdsERkGwIwVvW2EgvxzxZzBGqdUEfnM6tTS4nJTuZ2hiW6Ss3wh
z92Y31dcFOsTpVgkCTgjikZl330qUbyZjyIC2i4fjVtTofdFXTo4MVbHBvEzQY/xFt3dVlj7Dp4o
gIwUpS3HvRHRvvKo23iRfpgTN0RYVEghL6ctcJc4RBmzuZ2fUaFeeSg7hjpjylIXXZ9hgEHJvF8S
bOgNKP8OoQNacIZFakyrndlbMGhEYyvCqJ/QWoRZ+IrA29HWvm+Cw6I693WLM8MepuEPB1Z0dIeA
rtiW+YYlt6iRWwoqcDaO7r7S5FKM66t4FCv9Vrd6BQR4MEJRN+/bNPq93sIKafBaZF7rzLU5SVWu
J4+4rIbMvd+7kZSChQN+UodG66AVAakBkaXVsjLif87zLYzpPsGREXE6hhrqIuXTK9tE1j35wTCl
8AOt0AvcOxUSKfivr8uuA9TAIDlSf4zPCQPBOJkXgNRqkQMToRFBq+emlZnsPvkaigH0aC+U8LB1
HOmug75QlBZmxRhJZzY45QvvhnYyu6XHzzH9r526KfjHiAO3KoMAGf4eMrNKZnXwzhv42mZxCv+O
jRKKIocWWtosL156feDBMoRcwbhYDxwhz6Ro/xbK2k4JG4oKjm3u+yiEaYk7SN9SL+jJsbh3DusC
Y19Xw8C+2JvIRdyKoesyIW1KP8jy0Ar5sut1JKU3zcKOwJhL+crhc3ogZAmMd6Yd79hcrktQWyvX
5JS+VkZg6fxWWSMeNHWAtEmMdOfVvMKCAWSqjYSO6g8fkpo27ErzHrKuNvWTrXsgayKpIkYycHfQ
pK7RHoCTgbM07hXAxz24vlTtsqcRNsSED+jQhruNGvXcWA/uis42zAqfxcImOJm18cjxY79fom8c
awbTrGBOfy/vAURvwef2zOi0UoQvCgbY+7DkLOZsZahOGoOcc+S3AOz0Upz6xVy93arwnBsvJcM5
t6pntD09kPfRhJHHzAOuJZmKTNbq8dOxjqv+J1lDZL2ixCOFLMtuMf/So18nLmhc9o/tTdqAvoa+
zwk1X3LdQA1/LuMyqh4MkSpB9HaLS3nA8bIIBQKeW/2acofrP8UWCOCn7D2HeyWnzJK/myubfYWq
azSbdea1Kx6CqFmbqEOozMXe6xAbjdsiwg79I8qk6Z0BX8uBRNG2K3X0qnZ3j+e58Fgzvn7qUKMP
Ra8RPU2WOcMQdU5Ksp+pwZn+ZplYCGpAQL60YLdm1p5vBgne381nUFHvVmAr26Pq2HYu0neVvWqe
UoHYNuxlvR2LTDV1NEsqLyFpL9ZhgWa2zfajFmOXEMe4lfQNq535xU4DRjtBmydSCJp0qpo5g1ds
acKIxQe/YiQjw3S+xBQ6JeUu23ryJGKU2RxaJUuGr/glTd4LoHwpzUdPIDlsoek0IVJ7hcpq06v1
oVFmjx428DE5EZyt42ANqDe/pkxHK02y5dl4mp7dOv9AYmgUXvJv92sU9xXuqoIdp2Y1S9v5VWPJ
6rjp8t6EodRDN6esfSylsLJcbO6F18I/zFKnr7h572a7R0ALRo5ziSIJFBWJV6qIOB+85fUu9xUb
WVIfSS8PcK/FXwmTrTko/Bu3q1IU3NxSktWqnYWDEScwMAeNuo+QbwWvUnTB7Kl7MKhXzQqOAJpd
79aK1rmf/rxUKquzl1uXxFPfxov9A+VnPs2twz7VxdnBBp/JGcgQCdKtVpgr3vYQd4GVUsojWkTD
UyaURbqs+ZTUvT9Hkoz+Y2jFKKqM6w9ljbOsF7LWtLg0GboHrYGCus3QUscJNMt2xS0edA0B5s25
UELaYeZfHQlNITHUwYJNbTcn4RRH7Vh98B7Q2z5u/DngudvaInDmk7fhDMTsGpNhww2i2gIC0yrZ
VsniXKytZHRUABtD+QhzDRt9LiQX9jGvezz+iVewk05WJ9N5H8hlfeXq3Bx4QMxpK1Yms3vZMPCI
kq3FTfPU/M3KSsoXKRUeL6JeW4ZR7/4eZzyKgni7YrP0ANKZ1yaHgFeqJMeDnjeTtIF8MxLZm5ka
IT9AfSLZsB1QcigcADI9tMGtTMqY7ivP/CbV/FAtI3PiNvEn8Os/M8T5YS32lqXBsXwWZbyQavaQ
yOA3MIrFKuWzlUy6kw/rcUkg1fWaUBP9LzJSH3QkzK0/tTd0uUxaJUaZiNMNrMIqgLvd7nyfsJoZ
tgp6n/cs3zUqOR33VmSbIAhjzckqY28L9BbQMuiia6w65ZtlKbM8t0++VyqZbwV51jO/AC96Ng/u
MZqK1yOz486eQqi2gaG/rT+8ySDfvv1ya0/0GZhqLbDoTMavp4QTmxxi9gPM88y2kzMNQhr8f55y
7JZGc5BA69jk44NRWtwPL6NTeA6xojwpSWpL1atMrKb63U3KjEtghFc88rbdrwsSWvCE+Uxn6yvG
xxIn68FeDFBHLGBgEOiFS9WrftkQhkEPPNPVLitl6/qCbXeSE1+B/Pp6F1VODnIywr3/vG95X8HC
AgGp9r4X4y2rPdw0o4A9Zrbzpzcg1lwR2YgZ58yacaKg62QTehJ1zjWrjJ5SePlmKrKf0TG2Zz31
ujDS0SMrJ5fLcAkL3qDYmw3JTLsA6GtOHyb2Al1KfkriKz+n0oEmj1c2NskWD1ky1UxVXIVxB57o
hCOr8cQqjDCyCA7iQlT6bWRVWsHRYE11lVYVzOru/7JIJK7EaNMPL/5G/kIcvv0Nm1Qb0ljVxw46
VxC0thfSESU45QUcxcSFByB6X8Wo/7bENlGXjJLE6aZJ0NPiH1Qf05iZw0VwCdr9vL2pQvgWiW+4
6NJ3O/Q8NGPpnnYUR5dHFr6/vyrt3CGrR+z9APCqcNN/RPWyfeqU9GQkvFHbKiBj6DipY9Fgj8TF
xt27nyWIuVGrZ3KuIfL2SW1NIjte/4okKtgELP6AQgssquH0V+utUSdFfcZx+PoijF2YYTSvF26c
sTTBEo4pfh1kpM9CMUHthZIFNQEaxbq48aujF3+XCQ2+4TuQLhYqAc2sCM+kd8qbQwTuM9B0Ij55
igLwKjcS3W6imi3bRTQvHRGR72RTI5yfxUPRDgPl8CFp5vzasH7N8+LTPX99lo31TAVNBD+CUv5v
baSLuHSEQ/vfH99mbW5VPXXbkdRA1dZlWMHZpZpmd8ItZ9D+X0oX6fj3ofSXBd/YYQIARH/FRzcY
S/uufb2zbPp1rqL1FK2yHVVtRvBxY4vcE2FVjCjDPugtlL57AS4rQOGQnBffs04HHlg4eEygm8dv
hh+k1PSRobJOzSN+R8e0GADXR1hEn+yHe012g4AoEiStVfJMwcK8k6hhr8+N8qYyfwgmkOzKHDMf
iAzSyXsJnEQYcKF57RcymLo5GDUYJXj60HqVchlHyznea1fOrSHKb5a0jrhXQpfBImSnCNWysW/H
zcDfZUUjjKKmrZlOAEZP0Wddm/lELtBerDqW9fyzoRgSSIWSvzNcBU/Yi/2r9FJQe0B0G4lkBbGk
oclBQKnbRdR8ZQxXiB1YGBsM++LDpZdBhL4rncMS+NAJdxwsO449+q+q3uR7qQJXmC8w2yfQgucF
9QVY0tHigLZMOafpsJhLg29WZCyEhj+zJlyWvXti9pChA/Q/F/3rBWuUI0TeOqF5m6ujzPTEnwAK
ryhEKz19rgYtj+D2NZQim7iNkIz9b4CNsk3p14QOmzqp0O4PqPI3hrfCYkF3cDQAnNAzUUX/l+3J
YvUXW+BNC6zxtcBf5VGh86qegaVGl2f3PZQsCUJifyEy+ItnG7sGN4yENwXwGjEEpWPag7BA+ZQp
3BdTgYKe1slv5ztE3Dd2khjs9sHJW28RrCy6NYhvwrtRHThKHC4Tn9J4qwFWkKAUxHQCrqhJ/cNq
/MiiP3quGtJJQPVqh00RFbVWFYpSgH4OWscTFhzRjUxULKTugrXZVdDdq+lTAEnrOeHmmP+pbeww
NMWNKh3ja3CI/R3A/OgSRPVMywYMHmB6cL84e/SEYoiddlAwk4v6oQzMpnz8lIN278iUNf87Cyax
yLkoCCkU3/dEb3KmvDATh0jiMJ+Lv+IY0WXnt7kZ0A9Fbon6jjm4/ogB8NrCV4K8Njon292zrRnU
I3xiYoiIDdJ9I9n8XwQmF2s/em/zzWL8+nuXRDpfEEn7OafDYapQJbg1DBlOIWpJv95r+UNRVcxl
8k5/n122P5jwUQMVm69zSuy/GKxIj61kAvreCFF5IDLkLjgW0NjoBayyDkYK+6l/TMh67T3Sz7e8
qhFjhALundZQbMFQBWbNwuOiT+FIJxGkzKYma2j7xsC3W5BEvRgYpctNFLYhmSAFU/AN/3pkX1AQ
0vtyXTq0lqJJnW3T/GsEzvfvjkdbPAAgIFGpq6ckGsE7HqfySnUb3C8jd8dXOKaRh4WjNMjDwg+s
OnOvLYxbSPJXiqQPTPRo8f3YqNwSwekYmQdFI8h4OSJ3QI3npw1jbBe3OwDQ8YRR+Fcj68vUzVsK
FYO2rFo9zfMG0QUlVjmxlv2ZuiYXasc5LuH7gv+eDw9s15AV1IuzSonOjmNbn+S2c6z5zTsn+jbJ
bSRqO0NRiwshudz1jaOXCJ5/V0cU7bnk9tftGHyB46KMlncP1D226HVplht37TZLbXxLUYzbyp6g
A6n+CKTWBsQ0TxljOxBurti+NB80VirbMVV/iKFQVc2xMGOQzNOVfQ0dJ/9jIPrK4W3p7NDnRenB
D3Kb9pfkJs5gxUoDNPe399Ao9fJ3HviddVF47SKjHECIxtJmG5N2IiyyFz0kEs9T3KOhpNVeswuC
OULpLZXB3/Tu0acwUzERp2Dsj+RvzsnoEz5Ev9iGuOzd1xXC1xYJUGZ7OGi+7IMrJo1SFUjPH+TZ
JkwEbM3u8KKxYrsq8hl36Ointn0LqXUFdaiGSknRuSPTJKDZDQjVkiNuBO7qhKtPbXynnKvT9K9D
zNhAnmbwyfu6TKhsqOiz24hUngHLenQRCACPHGGyYhKEGmffJE4NK5cmFHsNJqDwyzycJG6cbLP6
xgDuiiSq0COkybs8B0ICqOL1xvePB4tzy3ciywh2GZ1clyxwcmPvVsCL62ZK+wzFIPtlNkUmGRev
O77l4vXjydPChZwnua5mS9uEdwwKaxnGTJ38ggsfWFekmO9bUsT0juU2PKLFike16XF35zWA7tGo
P+iJX8k1d323tNgM8YphZcdMbyrovro5JRiPqxnVRxJbwo0d86t/p1YlGkByftpWDBsf4LQJNmh1
ipS8PZcSLoBiHLs5Ehaa0Vrh/vNMrFrjAWMGL5joqYiIlK82Un4wbb4tCYApp0AIh9xUZLub8Sck
/BJ7q9+aMCOYMQ0r6feYdQ2c7T+o2lqGH0A5UqWPsgLXheRpw/nNOwecC3EgafbBU0SL6zey9P6l
bWM7rJ5c0ZjvEkbifAsx8cm2HDiuDWtBZCmWdH/wP0hHE3pvKoQs7s9HAnLLGHpoemba8jTq14Rd
up8Sc+om/nPagWOyp2EozPEnrPntM5lslmKqzKRnSzUX8eH4kfl3UqHFHfHLLfVh9hwVm938vqvJ
fSofR6tUGyAwDvz6oSYWaQnd92KFaBijPdadVcDYUlCmZQPQBz4re38adid7GtAIZSGOdtruof8O
PVrbBWAjsgduPwiwJN2N+MlpbfPrGO5yIbzNjNNEcjBx7Em0szKys4PD95VIVy4xlMirPXsPCqjg
62ZPGG7rLT+jZ3YNzxWJNgktSmYUnyU3J/n6FATzIcOzTmX7F5GJfNOBZ/W2g5xFxXxECtbWbJ9g
+DvaEcBQ/oIfx4tfCADjOWM8fL+3Rq7/wJFyu2zNFIvbnZ1nuddxmfE0p/xRaOmNp2awKezg5rPX
rRU8jYTur5yQbL60QQRem3I/JWcjQgqn/jrtPTGh9yV5Rs9KRCCCJU5zNhRQc644dfs58QjqPG1f
vjIVXrN8La9IarqvE7GEfAXSo4HGxOqcU6l6Ima571roX8AuImUZEF0Mau2o4FyCKciDfMAvg4AK
AJfRSsPbaVtFPQ/1PPCuxu4ijMEuI0lFwTsKKt9FJnYUdgNF7grmoREi74sM5Izh7V/qmQhgyzQa
zp005e8wJoWpJtr+d9ogrQgmLs4eJQVfZGAE78YwEOOimgFAjP1kA0IB4xj+bD8iQVcI07wz7o++
hiMR//yrIFgN5wQdWUwpluX6qrdsbY5oFuIiPyb6dEklKws3IIRtG9fozsLHd8WAFHn6VCKoqFU2
67sPC3EJtKt5hv7pfclgh1fSDB9dVhLoAB1uHWotg4wFeaY7Iyum9A9hiaR6p10rCS1ZPdKmcsbo
Eto8hEfvkknk1cYSkM0ewMkwIKk+z3nk5QOrg3+3H6Rd9gVy3KZuqlMXNDvH3O/Ri9SH6x82janZ
GecnARkVPrf42INsIPUQ/PFmf3brLHViiA15ygSWRw+3KTZ3RQxhNWKkEt215G9Ivj3+keCDBWmv
bEDJ6+udtqGYC2qRiNPWaL6/7RvLnOgnMs2QVUfQDpPbTL60Y1d41gtVuFLzN6NOYPqXBcmZCHdm
1udBq5enTzT1k25wP6pwDMdiM8vhM346ndFiQzV+qF9yEhvDlKoogEB4lxzes4jWhhOBuyJ5xX37
25gtZtdE+PIMCodym+7XjzIz9DXN6I3OVxMYFrsPMTdtq8TNzlFbxv9KxkuWbBus1Vj63wf0UQiV
Kl8A62H8DnHP9OsV7DdZhDcgCA+otdmgLZlYbyFNpbIo77r+f4xR+WK5ASg5jtSmoHmKjYodkVFh
iJx0+fGtZbI9CMooceJXauClf+Sy0ZeStOKzeYHDPtqDO0qD+EI86Q9Qu65kHaDIRJgIteIc9Tkk
MNE4dzTD+kD/q6hk5jcR0e2AXBzo8bbYlDr8+rZErozLInnDicHvZX3Rj9QR72un8b3gvNpD7M62
TbcDQxfFv8EWBKeMmhtoWxVZXhyPAKQgZwq89lMEXbleJNLKIzWz1WT5eQw26u90BSDINrUioudZ
BxX76nr8Y35/j2FdCZI2w5FBPoAJxKGWPtjBDzKSdtE+p95RPRYaDq2y+sC7LdhD1rSlSwchG4CW
jVeMBqsJrIqb36jJhg443XmcJPyF/eEOihEUYoDJ07LRDpbtsJ9fBh0751E1HXDdjh6QGo1gHwv0
G66iI5aEs37hoDvNO1Egc89soLIRyDJWv+htg6K017Xo9UvOkvvAFkhH9mraYd3PMcBrJRTYylGi
LNhW32GlELat/pWZvINBxDmjKPjK9Avoj9NAkAdumig0ZmiATejzNGQQkTTMF7xllSchK2pfTt0U
9uzoAnhgx9QSHXRms+GabWr4WD5HG9j0NCQsKxYdyxacKQDjjx2xtUe/OrU0o4ZxN6mYMDNsxI4k
2paMaZO3MZ+xHO6GbVWWi7SNF+MDJTImu72WEJT//Q4rDSXTjsP8sZldIM4l0j7y9/WJ+OMtrWEP
YoCETiO13NxZPFUSqBFY6szrhkacsYIUkwJE21Zwzvdt77DBDVXWN4vs0cqZo5kDweQAb3LI+66N
S8PaFx6uzPTYgwxxkyfMUxJXxdlp5WBLWXC7Vvuu+d5KHAh6HRfa7zs6Io3UKklPy1ZK/jkwwczw
55YgqLeQOM/+bvDmxkKBfXCkMFJxukBZeC33DbFirCLeqHzeEH947AuyoVVsHvKb3FzBniBLCAXx
YQBDklmabQFMN9kjRTxc31gnmk2RYK8NnX0rmN90UJ+5zl6gMCBYOM0BmW2VRzS727K6HFbCglvE
6Et6bhT+rZV5uZ0ei2PcfEdybIYXysJh/L1d28n8UYBfuQXIiUT1rsuitYPUDYmFDgguAHpRYv0t
C2V44HaXrM8msNcw1vNPWMnVImgO1sSVDpJLIlp59kx9G4fVcn5sqRM68pFZXfYJ7y9pMMU/8Uk4
7rd9M6Jpxq3aKlHbCWLvolPDeQ4nSiXmRgOeShK/xvXAxhm+ADP2W9RbmL3rTKvV+V4GmUx0xhCg
Fzyp0zj7QKRwsGwFbHnbRlk//gh4hwmypkOUryGwB01wiPzmrvxuI64cWpU18Ti89N5wmvP+ZDgx
A6cReZaIDWEaFxm5o+23NVy7HKaEPPBkRFrLtuhH3TeaK0U6KW/CjUDk/YGby7FxPQNqR1u6l6Lf
tjdpGyYit1KM4GcSfRmtT0YfCQwqQxY+uf5RVsGmtlrktaLsKOpHpYQLimE5vW9Tz7gI9T9uJg37
Mk/EcbmnyrLUEUatPOiyueEgttQAFbDZK0mA4pviDnqYakJJ96qyVUn+v1WzoSJq7+iNNDzYHU36
7VsQoJ8wAgZ8Xm0G7DSeeh/O//pNvtOdIZzQucLZqU/AknQypuSuLHcAZmmfcgCIUxDP0UCyFLeO
b5BHvO/cKWFvV+wBWmlsZd2J7Jm52/6ez0cmeGBDiIt0NPkkid/NK8FJIzPpnt8CVbMSJFQIMx0V
U5gQlZLcE+LOezyVBnxc2TPImqMgDnqy92L0boDNWmSGI13MiRaznOQUohjxRrKwWFCs/YaEYkpV
qQnAc2FkBQGVqvBoxBjxTwwA+bHGHjhtq/ofXJclx3YawdsH9lS8l1kjTU69+IneohsxWoG8CUbG
99PC6FVnVco/YXNbSmc85IPvdDBWtmxfVQht8Oph4djBWl+sHtZKINywnzCmYgPyLTtGw9MpVYfS
aUvn36OmvhxVamgy9rpONNuJq1sLu/8sWRb2gQ0QG8OepN+ADSZ/vIIaA8u3OVdTdU1eZ2BF4EHF
blN1+3TYYcig+VYB6YMh5NPYBoY88djOaMkhOBSy+9nuObFqLIuqi3qI9NjYWM1oBHlwMusrEY6k
inRkpTCco8SCg/+KNlZJRmoUkzjnAPN6LcfnO6cy7BwwWSOOxlMCmoJ1LxZy57d98I0zJX5nAS1+
Ik0ZVkeLGPzx8JdB9HtTc3XNeJsEv52JxyIO1cWfqKH4E3ewDb02A8glk0Wq/xzZSaAnz6f0QEh8
4j7NV7pB54OHf9aKPP8HkyVJuYFReAq4hcVpATILA7lMst+1VZlj/LvC6dxeHtLt7oUnYkfyqVgf
qNaYXOuQ7n44EbCUllkEC4IIdMLJaTMgsNpMBxWoMRHHHFRClwejr2FJRonnpM21HfvpQ62mb0Q8
Q3T9J9pHPPYSbB2Bw8LhF1ZoJSvCwrnJEofXK3nO2CZklUkVGqM+U5NyrvkXokTWGRSkZOpNACKO
2WymZu1b4Fb4WcgKmU1uU5Ag2Q3O8uI7/eA8JV7IDpXTdirE6NV0STppnCHnvsXiaIZDhEwMf5JS
IR3iT2kDZ9ldJx3lzwIg58ugbFJFDCOgLtlZERoLQpk3riijEBLqodlQNuUMvpBcEqcPYzFtxJm1
/jjl9vTM6+WCv7tqojVm7GyAKXqad9j18swMykF9KKAABlZZ4GQxpGFJCyfnnrYZsapgVPJln16i
2Wxkt0AtcmNd9D8aWYvapKphwCRdlRR1h28c7FukT1fV9A3Bs1wCQ+KVWTQHQziq4oDjd3ESyz6J
5KTIHAXp9PA+tZ15y7lEpd3Yo8f8jPm3c1hTF3cbdnhGU0C1sDZmFBBNL6lRmZQD3nvopi7qCYrf
D7tZ9v/2ywQrpVoKlsIJeDj1nWLS8e1UrIQYa3qSMH0rPIt1ypROjg3sdLl2X+23eS0pevEHMoRv
1i/hg9c77F7Ho+LTSS4NRlYqvlySGzkKkIy3bmsVcCjzj7QktzWmKblhNTLydxWCRWbiR+F5KzNv
9gn1wbb3dAU9AHGcWL1uj8qECwRtWruOfqBeANamX5oOmAvTBx3kZQ7W5uG9pQ3N23IZOtCKOFA7
GGa4EkbQ/0VQCZ5yOFwM/jCHu5fDxIaaH5sR7Gfm61I9p0yCHLRyGf+p6QjGuxOu62WGq7lTFk6b
JRkBz79P6cRZCFfT2qdH9ePM4fTXfOMoe2xENNk0rUoMLvak1v5hagYRjb7ip9yYRNM/mFLLC+fw
uJWP2UW94/8UEgi+iAiXZ/SKv2kQeHXWnLcgOuYhXs4dIWZN87LbIaZrG2mXMBwloOMPdGHaHCRb
5Eg09tQBlbW1SpKPR7VOO6eB4IdS86RWQe+ry5Wn5lFCJmFqaYwjtd6Gt/oWkTjYAaBoTghlZzVq
B4g1cw9C13u1bB7q76j26Xp0IQc+h9sgFvBlNFaSoCCKvh0iXwSXoyTtAWH1lPeXboFM5NV2rNX5
74f99s8mtTicREYCOq10G5G+Elv5pB9HQzRDbQLJLFAdxkoWaEAWtR6AH8O/MrZXI/IlXpxogshL
gf+Gi5I+aumlWkPdifmq0DUI5N6fDFhhl1l7Lrd6ddR7q4GiH5Ii8/CekrGMIwBSG/3y8QEIcxis
BaiO+pbMfFLgFY1KHUknqziomoCSYyWPUCZpNn2sEkS8XmqNVBxclAO4JLSBylzGZm47sCxJtTKR
lgqIOQ5J0Kmf0xluLD80TzpE6xkzoB8BJG7JTdR2/NPNtEe1WU3TdBjlbuLKFvH7bIZO0yjmsKnP
1LJQ6AOadvIXUP5Ffoi6EGmUpmLtegpWk3esEd+Vt5UFg1R7dAWSU4liLjHoXvUGpKlZFU4y8iAJ
luk4LhBW76au4qkStsqmrknfHqWO8hrwDKsH8pFSzXNTo2Fhn4flC5lBHGxD4awU1akVJUQaKes9
ewM3DxMscR86eCZ/LfBoKzkVdMbuI0AX4DznZcbL0+R53xWmwM/xTSe/r3PhWBRlJU95ezrF4esD
o1GLcgBXH6PuBnV04tLFjcNV6ZZebeM/c5uUnEH0tVfywEI0XDWC6/3hlqHEY2VqvH+aPXHb90Nq
g299/W21t/+mOgkIND29FEJIKem6zG3B+HUxHx7rhVtlP+15CZcyVT6JW2Y4JBOotQYQYTV4KGxA
GFTQK47SWzGiI/57cuAo6LG7oKBpXSmPp4+EvizuWjpwmBXda/LBKg94sB/QkL13zRtVlyr5Koab
EcLp87qKXqOft1BVelEO6tg+qA/jBc26euQqK+bKb02hP6pysUkTpAQvNoikIdN4ndfZHwHXN9hP
9a40drJbKZ2B/nA4sL42tK4uBUJlEo9EvOp7mNcO62QgPgGCY6z6pcwnsLm8h9TvaYLABcA4ouZA
b4qMVdCr07qejY4MbYzOBgBz/Nm85vpaC+TZpdMQHOZWxHxnqohxOuNipTjYh2YGHKVbGoaIaMl4
A/j30rWUUbfQOaz6+Mo25T1B1YyxqzPoEmJ+CcH+pp4DMVqMMwBjnk9FRGTxk49+RJaXj++zBNvw
Omk7Zs2mHKgayZKGIykHbDY8R+SuVO1RhGKGcohnQdlAxzPNYSkDmf+W+mZg2lvVzI9rSpHtFY1L
JOBdyAnkvfm815c8qWGtjhzWWgyW7ZcKXg0oyWHiY/9JpIbAz0zP/qVt0RhGq4GlJJS478v38psd
WpxAM9Jyv3CmIpTAzcD5ocxvsfu21Luuqg5OAIEhl8v1SdWYaUEFZ18mVpuwqdMO9XJGFl+lqxSz
pqs7m1tTnr/4fz7EXwc95XOzROEMkM3i6AOox661Yi66fFi6Xor2d9wnnz2pgGs0sb0QtBn+d4vh
UE2jDN1pc/ICzL8R8YLxPLCZnfkCipyvuELmgB4o3aXR4Fr1VY7HlX/PmCbzyV4bTJhbf6poABa+
nE6nr2GiU0y5ACtOvWOOJNyKeRPQFknQXp8PY9YtZpu3jKGsyLKzCbsGFFQTn3N2hLw0QbmpsYJ8
F1U2g3t6o2Gg2TAmILv+mG3FQlSPTkDzUGwOiq6sUXpYhOOyWyflcOr4Hicv2cwO4pdoGQCGxFAq
giyMpL7JZaRzE5sVEmoI9o3kP7ad01XpEh3irG/OXRy3HN5G+VuY9tJhNXrhTYMTHPfc2dU77Rsp
ku8KwB1fnocOOGKp2pkoB5gxlzz40DHn69xuBhISd60S1ZyatF7swRp+iJNO/zfI2kBwNJKgwy58
NipRM3tIUhcvkQOMmWelo/BpeGvFfIA0NqylCCCClXsZ3oUfeGY4HkC5khP+luKL2Jv+NN93xzVP
Wi14Fi9BobfIbKGu/Jt/nALwmku4hDv1iK5a0/EqafOjevd9YUuu68Ow1GtsYVQQ2STGMzRYv907
m3YfFET3w3/rXWJIK6wBW8bFIX9hl1GCs2g8Dn/Y/zZQg8VKYeKJ8ihF+JqAQOa9qbnJsTUmOvrt
vJOYWikmAWgGZEesGjgL7NO+52O8xdES2NTBYLhu9R8ZOg0KxVaa48TgRA2OPb+8xGcVM7mlI/Yn
UJmUBto97k3OCIUnr32VpApjhCxGHLfc1s6ga22JWXFqit/dxgI5eoshizN6OqU6aypq7AYFKx0C
wgIeVznGtZWDVhePMZ2s46qMc4oDxXBRuUAAnfI/LxB7GqaLYQBHMML9kYJViIpSGsgObQuBVx2I
dbZ9cWxO5WCMATGjkwyDpx3GkZ6E8wZnejQe8mX1sl5b2wq0+WMsyyHGWcC5NTqeG9TW5OspqHH1
F41wV+LpSIGAvW9+thkXxZxsF3EFq7GYRzR9xbZqnduCxiHIub/N3ulairehzTXwpaOxy9rhb2pb
+wCsBqEmSkZQf++l8lVQrouwBMs/qVPeO8p7vfw/DW+dUQq3lIsk38aF4JTr7/eevetC0kiXGgPm
afnZqQjnZWFZvKZ4VWqFCVX1TaYd2xMbnjqhp2SasxfESU3wZpfmM9F2w0zmyDIG9Jz/zq3IMzkw
HJ9xPfp2sS0y1wqunI2qjc2dCnkg2bBcJ44sKucrwqBV+86+VoE1zsjKj7fT/aaiG0Hu1Uyu+89+
oAFmD9VgY5i1XrXa0bZmUJrlmPLYbQbF8BjRXNNeqKuLJoTZ3AohL2hOS7SAku/P2Rb15fzXOA0a
Z5iKWHe3ddSe3R8tzCqQPjAGlmoBx2ru4QrxnvQ2kxXNWptv01ztnVSaF3CUQrQPPkNRN/+kDYKG
jQlALcPNgQ9XVKVHNBq33RlWrIEmZXcbdK+IwTYwnvb57m6APMchb8022ngkWs3YbzCSXow2+XfO
N3V/8NXQfOXEn+VBNvgK2LWQPMiGWFNW0vHmpDkSvBWNptc7QYFcrBxPsRrEOvdIw2vQbrjp0W9P
Fn3Qo3EHvd1aTT+ljDVvRKRJ7UUqV53DnoCNuMiYfbaAU6ueY4Hri9ZCqDENgF4Bj9hIkKdRa1sl
mHKU6HnIOpxZDddVcNydzjOWL5xdfZeBzizKR4F1xlaeYofC9zjiSRDX8LMdA/HXkW5ORkIXqjNI
ybIGDxJAEqJW563dOe0BsdKzfHf9hl4qiZ5nQNMZEfCClFLP8Zj3O2661tuFQ456suxpYY4aaZQy
Mm9xOnJRhoLfCu3arZKxpUpCzFwFsSV+O2a3U5CWHmWzutHbrgIdrrzGBskakaTqcFzHHK00gdVy
rS+iFKew8Qz3wnEpoZBBFaJaiKRSZM0OcJ0W03KpUj+k41xSCu2K73N6REQcSg2JS/Gv5Eodlngc
+zgeMctgX0Bk/b8iBHhCIRZtF9cDpT7Iy3P/18sSliHILOuSrDVUkyjnLhWOw4GQH7E7Eo+r8GbQ
EmnC8tFx993vmbdhHyHjHgBZv+WmEVOq+GmLfzV7diPHbzlhb6iPMljQPjDizw5iFCFAeEArGt9M
+yikdNfAirYQPNaBvaKM7KqFx9O8Ha/I6YkvbVrL4adxPLXjNiW1h6o3BcidWQPFw5GLkDmMFDLS
7yNeC7pJfHfrs977AKLjBOeZI7OZlah3ljeg4sl5R0n/yGPsDNXiJgAeP/dwy4R2yU7RfSVNhA1g
jweS91ir75e5ZmGQcKTtPlvz1kksrf/unkc4HqZLbv/zOEOp0NXvLTKB4SyFgxrjpzbKshRysAo7
w2PLQYAr+UqzTKydRhtyfjpyYAG1afzmgTzezPck7cMfezXkH1UV7c3Mv+h7NYQO8voeeD+g4GcL
4FZYBObsMrAs7dWL+ralr/QjyM/7rl8zpfo/cBcDbilgaYsPFh6ZUbF0G2p+11hVM2H/U22SMzRf
x6W+DAg6/6yF5wy1WYZ8Au6Z2r8nTYStq57In/CG+M5EWXLG2ybw6orTvij0RF2ktxNSAWASomvU
rUdgDKsuN1MEKdvHa+lFBCJiSpXLpxl+DT/5hm+j7iUISdNRi12//3YLBPGlX6L3jnL+XWP7j2gq
Aps6VeuI/AyNq06DAOG4gb1fHSNMmJYFaustaieqVJ1smqicV761UQR1GHiEFTLj8fNShFNIoPLn
v/ta02ZugHwt9jRuv1pagOaej/1+KrB/W3i1f9aTSmtJb4KVdRlQItYsqjsG72eJpzAiVLFNqMUK
WweWa7KaQhdfffVcztPH4aRKQkkApgwCk68MAq50ZxreB1/YLbB5NH0AzGXeczSss80CTDi5Jrzq
Q/oP1RelZE+L66HX5G9lI21pyJ+CqZZgpph8zF/pihaPYH86Z+CzpUHoTGN4Z8mqgYw+tGABTkey
qhPOVKyZemTdwYJshkrQwRt6xHPqqtgu/N399Brl0hjlj3qdaEkfKCemYcG4U07jKxnAeqjRnE4V
27p5j6F6ht6yMuRmkhM2rTXkXg+WlXKiZStIiKPLHIqYFxeHp21exmEPOKDPbgmlmBdYsnoW+6Z/
Dox7RsjmKIJIOQhbW/4WfeoxhsS+RyGrUQEruUGosjbTmNO46fzmxOWVZGG81dXyF2CtJKgjjqiX
/ct3bhPLBaNucBvUPZxkrLm1FqVQqHEVy87wOo344eNlETl6hSe/2/p7iT2Y10Xp6QMQBaQJn9Q9
DFXblmdEvU/2zaPoJujpx5xCDTht6vqDtLEZIJlZZzKmnRE0QxZvgR3CSMf1z4lFWVUPcAxyfmt1
CdcuUzVfAFBqo08/7sYMeinuI83hjlgB9yuzf5NNSFng0sOczdo/IAJk5xAjYhXP/XBFunhR9VZk
gQjj699PJY2eRfF7EjlcZqKAHYrA9R0MjnUH3t7+wyJPFGJ+vv4yaaclhj7nwwFiFZlNSG+RgPTD
XIfb219ZVXMIEGYlG+PTmuYsruXQIErbH79tef8SkNK7dbc+J+KvIA3xxuTP0PtQ5KQ5Y3dIhp+v
+oHVQS19P0dxmvFG6qMiPlTxsDulvTY9b7zvpcRcuefAFiXCSbjeAt8U04MLffUKjSBGMMlUF04A
kZg9Q72Kv0bB6soHCyEyBMj9e6ljsWt+03vgSbGAyzNJVBm/clmnQf0wL8oJCnFEfjJbvExxsJMq
LQlh4Mjuc7e+/DsD0fyP6mjXtRR9w16+XdlNFVBXyo+Orw+J87Q9j/suAe9LdIxPwI5EwEGW2n7W
RH3mqQ0utdMG0oLqa0HSGxHWsfBcFiBw2TVWZL7XugJ71ZwB12XtemPme4uZcXL9mBT5ix4CCHTJ
mCJOxRpQUC+EVNrbCD3XX4qHjwsTbhSUeOvcl5qO4CPc4hQdF1oTFRgZX6wo4mn8ywP96Gnfgn3P
TWbDOeaMmgG2vq/v3MGCTC3feVUAxq4wL5Al11M78/qUIv2Q7iIEYKE+mvbFmoCBBJGOv5HRgemF
mdGr5Dr0Kz4zbbpnu8QY/NPIJeWmbUPV7Rh/CLZkNW6vfSdwL183Vi7onpjwCuOJU5f8NxeCKYd+
2/+BH6rM58J9hqAidAJIMAIIh3AbWFnOXGfwRHeFT7gT98BatxrE3KwqRyw+Qh9zMNDzHdAg6AKB
L/69nSbCkbCBlR24ZQi46RPn5ea43N0IP+k6AAhcOGrhOOs0k91WZfHsiuD9z0zOgRTmUzXwfKFF
eBOYs4EXBv0WokridI7f7s+ZL0HsR/3kamsP0ytd/2iXOwibMK7u0y5Kl7eieH0H/w8wKORwlomt
yGI2xUYAIwO96bUCDpy1nXq4P0AZt2UGlci/iCmBUlglOWwAeBHSloo72V+36NuNuysTr5savk+b
PBvWBumdBvbvBNjqBw2C7wIRnxcJe9X4mT5B8LkXC/yN/uWXGGLficAGPYzMk/eFLTir5yAem47N
EWQV3QKFJguHRBSLZR4xJmIKbuOSKr32IjJbpE/4UOUO3ZF8sGjGSQ0r6NfPfTpPzEkNwR0Azvwz
VNxUhbwTp+s/55zWT5qMH7tuq/MyW7Sq+ZzyXMCjLpjuMWJ24MYLQtnA6q64VRT4rBQmM8PebbRc
50qn2p3cXUn/m1MD/t+QaagDOu56x8EC8ATTtf/T+wR87+Y4qKwCI41Ze/Bp/LLlf8Su4pYJkqLC
WP/dfiv01TB8OYr1iYbo9R54e14LkmeGpciz7rxlaIeRlTiLkXHJWWA4+gmRv8Yv1z9DWpvXZcc1
Iobi8/pLIDYDSyOIEGNqEnTL0h/AJTWqu0Mb2vmXykSHRVa7Vt10aeuwW7VF9a8PsKyjadQAd9RJ
lYh9oYoAXQo7GjYs2bFaMbai7PYgzqkR2UT7ZGN0oXBvmsVNf9kY0Xyx3Ou+9zio1zUh9/wXxvWl
nfgINq6I8w88S1Xj4E3YBEDVXFo+Je4j8v8QFk5h4N9ScvVYIq0iFFGD7mVACNkF5ia/yFtCDti8
ea7cpLHOO6uXSBlFuk71gcwe5G5/Hgmm9cbfePj23WzcVrK4mg9PNf/nV+0AdmPVX1/8CSlwgjx7
UsxSLQAxa5ZZBxa+X2wFDs6NSmGXSPn2b6FyNdl5zBGLFlYmbSvutWLC26f3hi70xpraah3usMWo
uF0ESPGjdmhi4I1glETj4EvP2l8er8P7K4D27Tro6S857oj82eZJ1rSB6g2A39Pz2HFGv2WUDilY
Ul/Dw4H5PNfTASiw5JAHstbVrRD1XxRdpAMtdwgATtOEct57jrB/uZ7kToLocTfn+skDLEgzcOh6
g2Q1vCQdyRXajQM1S8ORXe33BNW2vWhFfKpTPMTHIyTvoNe+yMD9TNTAX/jX/CyqmEJx9v3H5mh3
ZDSPqjtM1hWi1XEyqooxX842iYlZgewdVg6B9Ue0d2SUjhWvA4Hak0WGT+RDEgQcEMEapJfMq+23
7EnZU6CJRdutZu/gR7JYsm+QyCxRusZRpCCW5nNBC224VBODyBIYrtw/bej1TUHVvsPmSlmlHicX
rIuQVGZ/M0+BOcmFz1tCz97U7EmREnaUHFSDazsMW/kwA8/1CH/v7MqVJ/JdWCZNtb1bqBgkJv0R
U4VEt7bnQ6RDTH7El10JSa/Gr09Nf7jdQq3Up4JP6coAtRjYkKfW114PnQq9bm1W3mm752/NuZ7H
iWxxVmkYuuDCrkyQKwCzAgtLP8fg9rGm+mQHsEk0k5F9UroGqZLzN8/TGb4PX7PbLZP2Ny664b1L
8rcNlPhITQuKBqBtKQMLmMfjmhUCuTMUOQzt0KHssBYwlQ+KIJ+CwLdW2rHt0B4Q8uch/51bVcI5
t5EOXluSYiJ43aKOpEUjh1hHEB6FbWahjmnXCTFJuEJiT90hQq/eu0U0Fxw8hk5IvBo9pxijSE76
R55pLtefOtlf2rhp3ZcOLk6Ozyjl5q4FUX339P2vQcN7fsZBnL6yo2G6p61KnucDC6HH8dDEQFAC
5VOB0sQ0RYiRmfc2v+uVeqOjAqvlK794yynlRHXUrh07Fet4zEbRfNyT90sUKHygvjqYgjTo8MfI
rg+8uPad500cA41p89iTZhoUJZhlBv85RaFgDyLk+gdiDHc5e2I80HqbRV1DF6eSDWSHmeSlSYAC
l+PQiiHMfvHXEGEh/FjLIWSsiKPQfnhOjBjAG7+66flBlg37t08O35yz+i1IOt5OwHMa9FUilm1k
4k7QlN8IAYLI47omOcuo+83h0oZ307pmB88LA9Q+rUZIdn71Ll3PTlSiREdKuOeJzblAmRg5Lt1m
jB9ugpH3llugjuL/XCQ2XaWoWuMwCLH+oqo+aF150FuBScZ0xV3F9eRQVfQ+741sZvVKoxdxdV6t
FnDROF2FnR90ncf4ZnDqwin3/OoSjVD+FD36MJghlaSWWuU7l3sRqFIx4cwWmMthWWa0VVST8I1s
cgQWIf1eqOE7jTFZ3yOFnuORMFQHaUavQoSaVQeFkDytT9K2HvxokrqjG7xFrofs0ahDq01rFcPo
zTw/pkR8ewsAIQlPZ0wlT0UfICEjhJ8S2k2NqdM1bVkzyyCsDs6mXDi87nh8eXERVVVBeKNl8HpM
NTHNchw+jEgkxQZz1jFbfUoZP9utwsfqMkixPy2yi1oM/kFCtbufJcRqHL4+8sKt86njJNEdUGZi
+o24/e7807OrRKFmlGRqUKxuKQQfNxw/arxV73Zt6ZmlU0m4Wex5aS7WBv3pR26/zpcc8W5R7sJO
JBijhMwd/FIHYw5zanJZ5uTHu6JlbTvmEPVSlqXHLYxzXLL0GLcelHBrXVYEtXLWbWLiHWdWRwtC
8h0t7pI+L/cnVK+ZCBwrHAjcvBRPr4hVaBPO4cMdM3B+co+YfFgdQipeM0Tc1UFP9/prFbfBbzuY
DCP8QB+z/RP6QFxiuhbNfcIVN8SLbpdH+SgxzXeOYT41Ts3q+fWM3yFr7A+lQn2QZTdiP8Y4203X
mgpSAhEW4IR3cwv58tu/qvIpQMd/T85vpbvwWyHbicIOMcf7A+OUWUuiktm87CLJpCrBFfmA6OUk
63X/Ypku3BlAdWzf5V5QNny5f/1Zrq8PsEI9MISer4ratKaXGnvgBKKhLhOwN3aj09f1T/Ohvliw
nybjGCaPeyT8nlR1QVohLdSEgcRxoXhPobWa2WbSvklDxL7rqp42xZLkVulm9LBS1rIYiP2pviFP
t6fKYCgMTvWxRWmAofKTwsshy+BrKCZg9lyxHOe0p6rBmT7AKQ61DG3rLcKERCJf+faXkTqFdJRw
jYpUr+Um/reDlm7LF0xF2PVlrikBQUyPksx07GWbG/vrEJxUxGGtdMV43QudUGGI8qsUpd2/4/Rn
E3Bc51lYiMJoVdgRmzpqh3NJYo4QJ0aabRMB0j5Lbct7
`protect end_protected
