-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OcpnxJkAFL6AnLMvXrz52087TjvkpEFpCBLOiryVKEsOqKop4+771jHatvsOOan9fve9lStNEofi
P6sCxZAgEaRUdkXoJVh889frIeILnRH1n01oAZi3nb9L4HfwMLukCmVjn7wGJt2VbmVIlF8QOsXP
4Qk5hE5DanrGiiwT+bfGlfzsmZYkWodbBKVZuYAqJSnaj0aXSQqHiOkY/cbGmKZoS/Qosa4drJHw
Pgqg3MHd6GgD9lals/rRkz6g6G0aVDZoKKNgs86R5sEO2Lpdw8ft7HeubNHM8vIv6a/hELo+iOW7
wP0ridXWnYeeCHD6cx/gsjXtrllwhLpyWIYNpA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
UR+StX0N5RixSF162doCwdNrQGJj8LUM9ojIF/tZqQjCE4lzqkj759qoDZXC1tMb5i9/xRBa3Uh+
uTW7K38A/FMlRARg7HK/OVQtPro2Xb0dzd4ZHMspXGewgl4ur4dybRvsuY84lQwxKmifuvELKtVa
9hS4nUEFPdEfcg60ZpIKI+6iv6iGxCqTTVZF+P++7fyUnP22MW2pRFj4QbSUybSmwU5ykYuC6Ow+
fyuJ0L+HKo2RqP9dvyLQC+uJoDQQ02IuDgxDkSe9gohyLyGOA47gNOqCHmYsVmzuD9XpDW4oTnwh
VgBHXllMuHUvmvTRFKie+Jhbe9fFvaiDvbYyqJdDprAMo8ir/+kQaf+mOLMKWmdIQ2PH+KOzjnKO
NBvR/9HL82hsyZX9NTAPx3Ugh/bjZJ6YWQDwxKipqNqMXBE8Hg2KElbt46UHPxq2QMUPe2qc680U
t0Rf86hEAXNaHldDDipELFpZb8iHEhSV61WneWuvEW8XOZCEdguerwMOxbDASgeLf6j4V8tW6BRD
s+IQTj1QWuH+fD0ZnqTchg7wZPcuhVQHuNQNZjjL0jonHAofmac5GGY2GUyfLsROG/9p9wOV9U28
mSDv3l+asmyVB5fd1a+XcYTA3J45DJoPeZ8VdGHqjMUR5ikHxtjcC3kKtDbYjeDmPSyJLyeHownL
0V7+Sm2zB1JOPZ4Ls+RXck/LSa/BLi10Aq4coOFlkaTLzgmaG/qnwW4ySFwTTPENH7aZJtUNNIgi
5eui4zq1H8A2Ckj3eLI6V3AgAXXe60t8+FyitfVUN2uzwoCbZ6Uc6z3VnG8fZygKtXzIYRgegWZ/
MzGb3g9NHLfq83GLIMjtbNlDMtrx3FHCy8a5kYUbRG6cTvyybjJ4pVakJ5PPxSFOTNO3GgtZ10/h
o6RN/F4Qs9u56YhP+mdtREWoOhN4NwqXaXMAl0m8xU0Cq1soXYXV5IUOcMBcc9miqTQFzo6GIkcD
INFljdBvxOAhcjxx35Q5RP5LEoe9TiSvofbdGcjuuTuHgBg7K/nGY2chsfv+zkA+BwN46ti7Z3sz
+Y0Pe0oPggcxUb8V9Zh80lh1onOBAUkR2bvl2D96fFugpzGBZgCXvDF/1csCyhUVAkJuM1/FH7DH
gqkQM6r5cr9AVEuK4nNg+8KWXDHMdgpG9hi8f3AxZ8/kirDvFH1gs84mVMtpcYjOtSVpVheJlP+X
DV7fid7y99otYxmkqTBwUROApSQPx2jFVUAdPArIToMWKzzUWBf4KaksLHsegUiNqWWUk1qLbEYi
TtOdfsyhFBK5hkNFWRkec1XD6TW3GiPzwxq0lSaVeZYxT2dKbjmJBKUwr2WjsehyfiNvpqCHjgat
ZSlBlr0AKXkGD7L6SjBdHia1LIl7aWB2AeFHR8J+DU6bfwxjU5okWBi7ktl9ODUjvSdKhLH+4Vek
tRcr6kP3lVilABw32dH0dcrnfQzdyBeTKg8Wjdy8Aai5zZmPq8ryA7+pnpFgdDBVoUdZBGMEDCXW
HlGqFfWZEGT+k7oy8TNnP3JF7z+SW5/HVg6NeFfKIg7Ro9Y/ZrjZDtNnRkOxbcykUjdjYA6cei8G
yLaNYhwFJcyqKh9a0/Cyx3OTz3YJLjlQ8tPCrjK5uEt8+3gzAvLtFyRsfVpeCIi1IWeHCWYg6Equ
ltb1G4mqsz/cHQY2pYosj5r31aS3OhQXzz9hJCd48P9we827zvKZpBrymJsKkkgXHsDvw5+cqxiS
GRQOCdKrKsUkWyO3Od0JEwWcz9Ntv9VceHBWUuBNNKskEihJlLPOUgfCILjkf2HcWkczjPWVNtLs
cYb4x/HQvGY9hoqpL3mqa2b1nfV6vuv1klju3tWv7c/CQShVG7gRTWJBGNodm8vTnnxIRiJuKz47
q0UlYkICCFi6aEBsdAJbmmKG+mdkY5KY/rbgCepQZxIC3rhJ447p7q8LdtF1zriVf6TDNXQx7YsF
XlnDwt32zvFGBHMAORfCVlE6JvBjXKadW1u6c7K56gjFK2gPZWHeLBuaAduQHi3ENNPiBe0uZpSn
pn9iWvUYgke2BJXvfS+MSGHvsuOVptvblLC4wSbZK4u6oTxHSEfqmnDeDKziscblrkjHE7QYBkrY
rpO2KHZgTzzhtwrNwNCOIGKdrLHCT330uUHvNX96QGGF0+sE9+vr1BPfYdqxzhObEX0d6hsaDm1W
17yma95cChacy+A00nqDFAACs5QThYcdyPcFigWaCyj1ZvOqekxhrS1Tj1iy6zqxzNocX0RDtM57
D/PKx40F0V2MdsOzZu7UfKpP6Xiu8Kz9M0yQqp3KzWpcMWvsfnA+nz69c5KTXfHhRgDxHQpq7J3E
29zMSSmVkeCr8E5DoQeRwgdZ2moi4dV7Bt54Yo69msNF/HbA4MqTHWI44xLPNkF2eaB+yC3B0DpG
QucaDWhDz+YCEbIqMZVS61hsL75pZVIFxlxs7TOCjZeroRIHgOVCJH2otHDnmTM96KN5DVJ9JRQp
otHxJbCJR7/L6a1rzAkEUxNXXkdxGKFiqizgIyE1uF+nAvy/ffLYWQbJu4PNANJxaBQMDTwQsGri
n7ODEJJFxjtpIfQVI+8O94kA669eXmTjwRwSD80ei/hVU3eIa55gy+Erah/ohBz14d7fTFT2K8zE
Wsb2f97avCB2uDfNWX+xkdB5zHb8aakQGNR2REGlehkwFgE/EsY/QCm/x6VZ218sv73URzRuK6Ly
efY8GBZIBzipjGhbYXJzd0FDjeKLf88U2lz16s9qwfZIFIRtOS2c2f/X5yImO5NXfLhv0UbeFDDB
mRrxLi7gBlctnGWzqaIaH2MF6KHn0evipTnCTzfhRVAmhjLGb82snX4DyajKP8so9XLWzErqwUjq
UZS5Fx/oSxsPIRQHIKSaTPGMMDo0A5eFjZVJByRiHR7dS/tBO3GY4LXGvJ2rLMJnIje1tC2yPtOR
UOqR7DxlPFbUyTdwxUOviCGT6+eiB4QLOX3Y5Znvu2RzMfnT+VVZUcG9sZlJo13kusx58d634TJB
hVwjmPgvAvRU6sgcaQ86gme8Fezl+lFIBYLKdKQNlALfv/7bf9M1VxWiYm7Y3VJjWJNpcTfwf5a/
giBSylb4Z7JbOAO3xRFG/7cx/oH4EdNGAl+Oj704xB3kb83nunJc3dTDthyo5gLZWquB0NesRusL
dt1JhCzdOL1r0gAvYwYohWOnYMmxzLkUbW4o0nKtoqc53wcnBDLjy01HDDWqysiYHTu3tX+GJSzD
VJIvXtF2uOTADAgbrY8SWKabpsfd+hoiHrQP1oRg7SrPLZyOGgE00iGcUit3TMaiNoLzhxTNqbaf
qaEY2qXEU+LkIWS/i3hHh/CU7HFf7uq+RnPoSebFON/rczGYI72DvLI6bEKN54BuilbXRqY0Rofk
WtNmYJbgwscZFd3QeE3BK4r3I3YDShpoul6J2PUnRkHgfIu0NcLANbCqoNLV62fqlzImFS1upnru
FA+oQkoUk6EYcSH/BiQbknS7OEBmHJO1mq/mcmdl+Y831/yBHDNywEzNW0nywpA9p+ZBTsropU+6
CFnDv2gUDprVCRY5OaHkBuZO3l8B7PrVvc5UTxUltFs0nrSF6ZDtibnwjt/bslThVTzCG650k7Jw
jAiySPan+wcFDUV1E/cgBuk9zjEUYwjSz8MzFwAdK2XdqAjnDEiflcB39PDcefDnZg1xAgg0JeTN
Hx8Xy05ww6YRvIixwLRpaL3cXyUG7Q417ayJnTCpFlXYQmWWoXRkjF0DQE5XDIN5H87vuUZtY5rF
Zd0FzgQow4I1virJoAzOoyxttGdAxy88pj9I4Oemw2YP3NPxZRPMFFEPXTjCqnMXWla56m4qlUq8
kUZbnhBzZoqj8YSkh5f1WAnmnYc8cFkwXeY/+lhx6u2GHaPltlyxj5oLGUM/FQvlFbta92LM0AOi
A9n3kBoLIjrHOFdzMcAll1zylXlrdJyz7qLAELqj4RACPeqNR+pAC6kEKW6K2KoOWcQY51h6ydA5
t0EgkTQeuVoydR3A7L2W924SEEfSlMfrDuvn1+FGwrTOz1kagwynsdQO9M1olCQEKQDvlGS70rXT
eIjboIMIeLbFXhsSD/tUA/9WEyb4eEOd+N9w/nUMVCcz3R26e/jOkWtZTGNnoD4A806ZZtefdUAA
YDrk+liP9vSMUpsrA6YKMOvzhY9lP80SfUFyDaoDCZA+qmtUbXVGokFeAMru1Dnj1a76gQCrq9ae
LEHs9Frx9sBs4HhCkE5ERI9zlQ0FjnYXfgvtCW71jrmS40itmfDCGy/iJGuTZIQNtI2oKsLZlMWv
bhxbhf5Hwx1SL/RZDJ6pN3JN25xMlqHGlg3j7VHs5nbl2VfGyt+0Q8e/5BokWlo/QQsWmjKgAeaN
QYmTyoojD9vJFnCMc/QyNbpl+0oWCmwWSltTCA/2jMfoI9Fg6sZPJTMIzgaWfVelOK7Tqj0cTIsZ
6qc5FrlS7G0AGPixgByoB8S/MislR9Y3PBtYSgzQtBzQH/y245oELAo1SUYVAY1+AS35D32k5Yc9
mBprQ+Fd5CVeZHWEoYqdG46f1ksumQ0L9UjkJBWD7H9rN9GeaXHuf6aJGrtK3gfeK/dEg/m4NjgH
+Gl76BtCcsfYl29IHPoL4lsPYrHKbLaQtayboarfCiPCJNZ/5xIElnII3/CU6x+jGyRy65f7OumA
2IBP2YF0nUYHhAUzNCUblUTLRtJxCf8ZCVlRtSRx2DGuFqJ0LxruiP5I8VuIxtW6YCOibZZprhW5
+hIQdi08l50yeRHxDVSkdqDqietAXRy3ryqMHgnasMab3UN5vcJvolkjXkKajrbOjVCHcA3he95F
5V7jCR8lNgLoi7Wk0O1oWX9xzH2cEdsWb6pzKOAmHkpIAxS1fu3Zn6FzdmiylM85gQmJXklHVqyW
XEcWyyv2eqWhtAHCfBGIrDSFJs6XnxDcW8M/BAuk2jFUunkUGHozBoK1cbeWidLFuRrxDS9H3qGf
Rl+nufK+e2OjA9677L1R9YkVB2t2+N1fYq6dCeXc/+1yOvQCwITT7+69oMYDK5sdRUhoTupUjpa7
f55UdZ365JQfUHZjuE4K7BPctZ1gNVvkRpDzLPHyF9pEBMkd3o2M/If5sv2ZT5/cqTui1Z/LSDoE
2Ybr4mGQ2rOK3mRh+qEN1di65miL4N1dTkuAzXUgQn2rEM1ITqApfdz1nk+uoKWT489QK6rbaOt1
KERwaPFcJszHjoj5yOEAx6VfHq7WNvbkCfAIUlrGTPHkVjOmc2SoY6KqWD68Eg8F2JsUDPzSlwX5
0b9GMnLPFKtAm8VW2kA8h112xLSaBfz/UnEi/fSuRrYHchj1TuEVWdzE3Ga6vfrHAlHM/P1/+113
5S4VCsRrxZaegxAMCIUNZZWZY9SbFRWa1TB9kQq3RPGFD0yIBnFRO61Xe56Uazo4R6knl8C0FXMP
K1xmAssurVgon87/w9BWRK22JPPrH6w/GndvapGo4mED4Bp4KjKsJT2K/AoXUaCsb+f4bBJdGCJQ
uPULNhUvQywwV3SSK46gLAcHaXvkmZcn6mfHMoUKoKLaV7Ov007NztusLMSuBe/22Y9oLofOQya4
AgQb8BP73Tq2ruoavUiazAvC/SGfh5wJgYHXxxSJXzdli1FrV9M3OJYNEimZLN/+RioLqYuCh8xr
QnmtMlE96siu2Vdz7Q==
`protect end_protected
