-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bSCACgB8mwIlxiKPChLmQCh1FATOIvsBUDXiLAEBTcKBsQ3VXLakjGt1/EIOi+GtXrMYBjvKy1dQ
HBiNowMwMja9/rT0WE571qDQaihWD2Zy8Jr3az09tcjMEoLLFssCKvJNcgutZDKg54EYQhoPbqmO
JHrynODhmVt+JX4Mspp8SJM1OtDzyiioJaA5XwIjKeYvMgYDDyhlYkHUn3xNdZJ5UV7viPE/SNgm
4EL8aQYJ1LQr9aq7Ya/dPbtm67jraTpa/mGIAMZSnRd6c0C1wpf+Ynog+3xZ5ugG47h3H22KG1ea
iiZlS1JCGaMolVtJoaq6WKvTC+ylBjOHyVkzGQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
cfzJ4qes6jckJCnvTyjjbr9z4rGbCP+eVchAcEaCkxOjYRu/dp+PxDVlZyqxUANaQTqVYG2Yl2uX
Xp2d0Bsz8T30JOMJGCZlwFxjfQOE8Rslp6w977ThDmTG1qzR6Imyrj/RayZ7YFJMMzX4D9dBqXZw
cjHetKkZDt6EkE/BQGFTP1WOfgJ9GTfSyA4+4VHHTVdi4Yu21wqK4zrrYyvW/XUbUoqLfPmGxi1Z
nMiyuIn+S31wrdkAPhwlruuAUyp1SKaZUsK50agunRz2Xbgrs13/rCyVY8g0DHb9UvbsWLpae7JT
FxXw63Vcn3LG9uji7Yn+3ssUSNhErm3icoRcacHF2zWcYMjJpjyC68HTtoY41Ac81/ArSYttozd0
Vkxj1VhITxQJSl3z3T4WnETM5veOw6TmR5+/9i4z1ZicVsWzqJj7jQ3J7/8k0KZ7xJJkTlaQEkFE
nfIyNQbTGsPWCl/cCFStN6e2G0l1d2sR3nLzgg2KpXkJvlgJp/VqrJFwiW2wZ4X6k+p9YKqxveqW
WU6YQMO0XrWyj5iJwtVemB10qYO341n0fjTETcIVBpbfWPKxI3mxxUWIhPF1g/VbXlIL3RdyxTjF
hA74bUOciJ3ZQnBssT7s3mrPSoei2kt+Qg8/1qx6JM9v95ISkBgSR6Q/vFU6dCpx/3GB3ye71xsK
faPFWDXYx19vqrjxTN8Si+nWlWgNoVdLFtuqc4gs9+nFxdHts7+o+VVsa8Hj5NDzA40lVdwxDG6d
pK7OMkSs9G1Js0mBqLjs0EXwlprOoitwsR9f6zWrr+9M5WvO56oroZcdho6y+oCsWPkT2ZpcsdLJ
f5FuZpnZEKrpvzwUfwCIkhmUEfcfanGKbkMNGMgpoOmI1FtJIG7ksvlbtHfIFD1qej09y4CFRxFS
bkpdRuAVlPPUdHdhqXtuN/Cv8YdYB3uabSQIZeqh1NmDz+0PmRvEEJSRWp0YPeHAeJ3dPAK4pW5r
r7IgEct5eP96hXkHRdgMyU5TI9DySVKL6Le+se3gE1yC795Pf4djqjsoozSpfYmVHlz9/mHA1n8S
FzBdzGwXoMfwDnsFsyeKBAtk+/7PM5T2i/agHxhPWPiMNUwmypV+6SkOp3f855dVupuXfVOLGMJF
edEaiZXwsJffzx2c/FiY4FADMIo58Qnl8L0yXdjlzR1KKhkHKOuMbzsUbTy2/31sLA7K+/26Uh6C
A2bTLHWOKlxmavUYksrKN7SYCEtU0dnTRRVmuViKVN3wiICxxJdr7me8qAB2L7tCXpcd72RQ+4YK
k5hYvo/T/dMJK6ZQA4twh/8XPUXAJnyQHJs0tFdC4SEioGMbHGgCnuKwfggoGF8ph9VCODJvRNpl
1PSmErNs/0avD8eiWkHkZYgvjvlYAfD7KnkK//lKdj3X59UM//Pm0XSlNKl1jGWzvgtq/kdAjOyg
35jknA1bVuxBy1CBr1lTAcZefaIjNj0ugufOfYz2Nkgh9j+SbM2uUJBdr06hAR/s8BLL/Ho/tu27
pJis/G4hZ/SPwoABxOks5EUt0jDLTbUdfN5rghZQTgV8QSM8lqOXbvmiMX+jpOiwNI7AM3KyKDpf
fr+VwE7/V/oXBg88nhDpl3H99dSQu3McbU22aGCC4vwFEAhicM2qwAX7ryWJc6LgsjyMJrpKLCTg
UDGaTKEvhrNMfVMlFMeLXR/VOwRc36sbHaWX6tRtbahrR1DPENAlJ2wu0WV8iUkHM/kcLGylAfvG
zDB8GiR8c5wbD51VsWdBUG/qFItnlnXWFqZKL792gCnjFtLS+7B7kYjbPkFCPzsyHoYz1AQi1sNk
HJWBYjDC+n5440hD+sbbM7uaxiujuPQtKCiOdYE7p/OyQ5aQa2gaP3PMifuSpj8+9xiNkHFrUZay
Rh8Rv8+/3XuVNObKR+3eFD9CLsVREoh/VEwcg4tnDwop3RVRVhYdi57TqjNDXxlpOZ12mePkmBn0
y1+n39GHTomqTATzh8kG3pFMIbR1jikghjiYXLPTkmw3BsVxH1aaVlmFNQfYOiJqMiqR0zqwUaYf
cqps7J30g3bez6W0GT8mlTYLY1wIHcS3WucneuKveW/PZavJ+YJ5eCWg1CkiHeJgYyDvGgauxWk3
vyO02cZwxuvsKIXo0h0iSqXvmCHzUaG8jfB05bODvZ8me3ignr6kxiiZy8C2ue7zzxIU3sHZ3MnU
pGBZjeTGLo3brVyzRFMETEr31p5NrkyeJGT8SFzhXl06IfYOnAs73fw99wpKXKVlsrzR1DxABd50
pZqkI7ZpVkNMen1wUyScsnltX4QSAFwbWxm/WfNqcILdX7PuTUiODOdBFJXyc+gs+yZcMwGLwDSI
ge8cq4MefPKDVylA+dvGuCmPdAQ3J7775xlsMARhDfVIjGdab+xao7tUrz1ePqdxg7rl5w8IBUqV
gRqGx7FiIRMR+3bd0/hCgrZhQjKLrfBOtaiEWl9nn5Y0jzST4JL9Ym3r33F15boufoX3diERIZ4l
1UgczAgOXf9pP523Ye6G7IdPNBnwp2q2a+S5fUssHFvCWsvY4pK6dsYxS7Kv3JO0SNXaa33LSYBq
p9zj7MRvyvUIqVSt4qk9PFZ1kz076PdUjTtI6SSsCLK7eah49pnueQriQ4BUf/ZJfFDLPVkaQKC4
ssxYzAV5OuEF5c+FpaFJc3J8pedIRcNnOPj3c6TR5fEl6ubc6UhOt8h4d7tGoNMb2fQ1aoz4HXoa
hiOHsEE9sThZC80J7yLcSD8mslki7LUr0MMBGvwLwmYIDw/T+XAmaX2a1pgANXDgD7h+2nNeIsGh
rsSvQnKK8tjW9v3FDkQs/slJAgtd33VNkxYbu6auChvh8SVbeWH3PfyxioSuEmotarKenq0NE/9p
TR2vv6L45n0YEU+j+6EpZQ7sRjA16T4ZPMBOmbdE7DYbsZVqr86tiAZ6hR5gm6vjm6YWFgJDExYL
8mWyWIyKAE6dLDSmDKS2SBVYEX7QlLEkAJB4DPKaRBVdNqt3Jequm5+YUToFQmsl9bacxYZoPWHX
VBOk44ARSzarT2Olvg1Dkrw++lfARBJVmAe6F58Vq1JP2xi1CGbENNSSmt1cCt9Oj1bVOg2g1lce
q+lB45J7D37keJwrNwr9YYU74SGdXeXe1mfFSKuw2PfZYuilqCZ3MTJrbFCSFgNXUIej126xPgSt
h9uwFzv8+Qlg/IvpOXQ0i4dKRI9rF7DtFs9HC4HsyST9aCYhYCZegPbumM7cXshB/ivFmw25Ctam
FTa3vMoG4YHD2ZThOEYOVjAOFv/adUC5eotT2d8OYf01+JtKbIyQnKKTi0fjTVdqGJ61Ki1VfbIS
EJrX1c+cBukoQmKXLTc56kG+wDBDlW7y2oG6Z+9NclGIOaAjdzVHKFuvGqMnz6bp29Y1MqesU48f
Oa4YpuilTGO7iu+Ez70aQRGOqOKCajjlQAa67a3PnAplb//7/Y1mwwU+2d37IsjHQVI9XxP+ltXj
MQPCrooIyM/GwSxKU1SEsFPlrgf6d5EM46B+UYSjFZv4TdBi4xpNDEv7bJ4Z4Sbaf4Rx7moA2HP+
ZtVysUWrnNkvxzS9gZhvTVJttpRXMZi2/dMPCG3GLO5D9E/U+xBKp24V3ENNScjBitIGf0LEc3ef
ZTH7e2FOz2Gdz7z2wWooiP+oaFsCK9bKxkOhcWkC7sNTXEZESkr4MUAf+xQHuiJnFYTS8kcAhCsr
TCBgbC+NpAE5O5xOIWux7OnmxJehXqAMzXzj5lv3ddSblEmk+fl1deUB4HJj213C//m+VAt7pNXx
L36A2hM+vXJo+83bmVY41jtVpbALTi8H3xhYZGp323zGsDz/aSMx2AhWODdFxJyHbGfzYC/fkSKT
7vHjW5D/cFmBC1ZahvrtFUqWI9BLxzCTkstCGNaXJ0JtVqMIR0M3qIXEPCZq4vAFOhIVaXADVv/B
QSMZVbxT7EUx25AOBf2dySZIyI4FE9mmQFHR73Mm2aYdsGa0P8X8ROBL/2PvdLSHpoqjne9FoqXX
fz0rWuM0xjJAhnTqUe+4cf32adPlhDO7nw4HAvmbtOaDFkMIOa2/Wezv5DMYeLe3qw03UJbHP/vc
lnAy+Up461viVrt6+8FGdhWa2Y5oeyj5Bprg756EqPxM4/bqR6hSFtCoX1TKsndYlgzp5BJGGcwP
G9E+J9FR1pfjZF4aQ322ZMhLLuoniqjGbVoDcMiFCgzz8uQCJZ797lJZK2j8yd/fqUBgazMmSY8q
s/OW047PVI9+IsRldV+wqvnWZXpwJFYZLGhWoJcKujQ88OH3/iKCyvZd/ad2gfCC5hksNPqKW+81
WfzlhzJlFealrrw6EiQHUD48ouQfMX7jdH43Z0Wjgve9wkM2/1GUmwtevNWr6FY/BVg6Cckae1uY
pvprKEClfv5fKGt48M/feelocU6leNHFb46VzRi+orM9RRlE8v9Lfa8ddksxrqUz30nApqB3sIjv
jI/IXIIU8z+x2c+znKSYlakSBB9Cl24knAm8yydccD+HvIOtT2WHLheAjduMzTqIo7NTjuTPw4iT
bLFAeZQZbe1+n4AQcoc632Ylol9M9Bgas0XuJtv4NQog7YcutRpUG+M+sQWgFQcTDXJo+S38OGfj
fnxVd27IJ1/wRio7YG2m4mFfyYWjeC//hRP8H1tmpAw66Ce7oMYPmf5jsxD7njQls6/VqctJ9sp7
RvbvEgHQa9sGfPCVIOaPHgjRojL5LtZ00+/E55lw+OBFViBM/DZwqNJlueIzl7WF1OpvE4uwZW7/
uYpLOM/HfURAwPnu4GQtLFaQhUqfI8ye4/mXqHQIbHJ/ZkaE4GcsXhIoqMFPf5vqe9W2erhSLZzl
FnysgLqPwSe/AmfZ7Igev5watwSbGDb28csf3i7Jx/Kx8040Hy0YVms8Bg+SlyjiE1Ou0QSJl4cf
wx7s9WQ8ARjCKsIxpKUAQbx7JBzxBLfT/liPpJLVLK2IqScbA9bW26S8m9g3Z6g3rfUv0AbC7QO9
kCKRr7h3qHpUbKBL5qGiTIodqDi1mPI40Iby1ZB59M9f3JF4D2rELpnMMhtsw/Yb82mMiL0Fgokm
gW04M3lBtxLuWWytB3uGMd6FcHz/4vQOFN9iWumLOkpKBMnKc1u9BBjXINRT/Is89e0SJhI6iotX
w5amCW7/qV+upruCmVr4nOSoJkq5Up1A0CLyDiJoSkYTvwneIclQgaPHL4XaeGNHDny05evv8Nm9
j7WaaGUPPBlkFMUCl+w9+cW/qyC0HE+PJ8TGfqHTMa23ITK7SN2ImDzv4yOZXCogYRo7bsRqpJPr
4BBlrtITmU88rD2yctW0C/ghBfVhhQfPNj54yGehU0t+RxXKsOyGPBMKD1nWCb9KZLqiZQjUHSXL
gytIzEhWqkIWMb3nfraQkRMeY55Yk1G8nk7KZieuOGUrJltFmtMCVrsGQXT6wV0e8bLEGbeSQSv7
hgMbrQlFnaQfBvzSyPk36ZLNUE2ZcOH5svMC9Y8i8LTrgtmMM/pJ2Ot2AcCQkwaTgJ0NHj3vA6sO
5Suz4Yfv5sYeP/rgvoKherhRnZR99th8EPcXEH406V2w2Nynx7EZR+bj31Z5XxvRf3Rj21iVjHXz
uyxoCMqH7Rf6y2/I0cumfIlfwTrsGk85a8aF+RADFfAT3BIfsNvaJqTSMG1MftZsfTIJ4AFxBO/n
U5974Lood5SJifMemDD0zgVZSXV5dsRan+QIyMKVGQVAVvxR7o0mST6xaQtjDXtZKgQj0RTFQ5gx
1+vy7B4LWyhzlczW8ItIfn8NUPaXT87xuP2VTwapJSZD55jYkcHUP4s/PG4VzFKYxVCW2ZVvE7Mr
Ztnv76V3FlG7ncomJoorCYVEHXozxLER/N9/tuN4KLHN4VhB0IbYRbDxmb5ZB1vbzj/6uOBLb+9U
Pnlk7zGYxdsccM4kcqkQgUG5mVvHl35WaW50ZQLIWjvWqJgAZj5ht0/LXbMCS6ZPTicFCVl1yFk9
avxKOGbSfKm9qaoPc/XLYWEHOre8EI8vyCFIIS+DMrgkszPINp0L8plkFcEjzgApc+3VGe4xu0Q1
qCYj2qSONnaJdWRQLkooqoNPPJwYaZEjhWZlLwVixfdO9Q60bKP9F4alrv4HQpz2L7FAQQstuj/E
xlQmn7Df8I2osxzNnEGuUmWwoPqBJVT6WQ3hMuYR18NTcfrAbF0IShF/mNW6wLS3xYZXgMjw7OrY
+LdOi/TIN/6BwKllU0xZCl6oBKEOh8LxfXLJSkguHWAbZumN1q5Avtsr/Iyzr+xNcMkoSVlflOSU
k6h0/vTPLwor7O6ByGW8HjLomhDZuqDjrAehdsvKXigelEjwnpZpB2o1oep7+hWtp9mOqfeTu1Ff
gWb9E+Ei6SDcnVl6KAyDzw6Ru63oui429jOBW5U7Wl7eqDiC82UkxCLYGUlZcg5OFQixvBHqxmxY
0kO6oms3qHJpIjdSXCrUsKI4BvKkfFSkLhSHE/s/KGVC46RK6hQweDgmqyqkwiak4NLH0fmhX+NZ
Jp3S2l6BeSCJNiy415UAw/qhVglJr5tuVBQtlmuozBneGmOn6E6vr/JSkpjWeyYPqlOqFnfZMsr4
UMkxwsfSedqaDZYtMNIBcCQL2ULoice2rDyG4cjzl8mZykCHBXf4J2ZMDEsQ4i/8AyMhh8CnSAIa
3gH3j6o+grwObBycgXeiC7nefG8UujiSPicmWcs/r9QQNT1JPqatrSuObfAcoJFcU0RI3uXKKwEW
u01GGBQR56PjwQZWcxDf/F+yWNLAWwicAQaiWpMvAqt6UYvoYgtaUpRwqTAdBWjYjEO8egNqR8tm
3Wmwq9QFRrTPnjV0cmy2Dg9nCKe4IsZUEWZ6ByMAn5FHhn4xxaf19N2/DZaocRHAPBk9aZ+Ghl/Z
rEHPShfQWR+qTJvqOhfrTvXoSca6l/TAU09zciVzdFFAfIMzkDVE64nI/LY06b1xypvIMYBStoVB
ooUYS6P3WdMoh0FMVirxwoKPzpHH4/tJey0+LIt87m5pv6jxxQx/0Rl9ef1f2Gndr6QylZbai/vR
HtWWS7ALLgNiRk7cSekMzab+cgiAWvJpcaTbYmpoWeYFwJ/dFc67H1+Z2RVoYuWZENwy/tTXeyqg
oy0aZfYYsqXL5ddD8BML7HK9QHZlsDs9bSz8aDHinVdjIrh3zSwo47oEOOOD8/EAbxDC2GHgr9mp
bY95VWkkE5bWWw4D4piHi3/mpozDl5ckMEwcF5hLF+itfRVuveo1R5s5rATBZ2q3HzXxLOElopg7
ClK8qr1A+6bNLRGgOuX1Z0+1mRf6URq8lDsyUPMITI3JWyRrapwxo3/g9UNsrLK6PWFLueyfes7G
k+nA4SUzmj8CGfJP8e1JObCjwOK6Hj0epRJXvIhQrJht9cj748/tfRD7V8S9x2i2lwTiyjVv7Smx
xm6Tgm6llWC/3vhEYe0Yew9LUnxaac08o9Q/Y7CuNbUt5QpN1BjW8qY+NOjdb55BntaGq70larTh
UKfYksm1du5xB7oMtWyXMiniBPuERvsssGLzYfkgnIpGwDxVEYofrC/bdlcEJh676d35NA9bXwgg
THqEmXRbcn/BOCVx/2OcXl402knkA9w352Nc/xc9Lr0BSFaQ+Ej3uGD6iTIjmUtZY/OsSfWnOf0y
AixNhdTb+mUFqb7Eiz5gL6VaTZmgV+/ZHJpSOAgaFX9BZ3l/UQ/RAzlUQaR/G4ztTTgS6hbXQdLE
iM/VYdYQ3uYN2BD69rTajphKAiCA1nxDMaDhBz8wttgshHQkW5Hq45BwK1btAczSkce4sUnF7+WC
Wb+O63oQoRVG4zdTXCMt2ZklpYJ7zID8UE7Qqls8PSQVl7ThAYqcX6eqFVVpEgNWHFh1JIWVHaN1
StQluqCQJRD1N4jt/qqOSHX8s7QQeck/KGkMeEH+4E50rBpJzMZ24GgtzNEwT9MSTBJaayNtV5+U
mHZd9VWc30Ilx20tgKydzdW4S0n9B+Jg7QoHqpokJr+VXh+ePsdBwfkeEF4h4cGSzv/lmz8kMgF+
bW1+8tK7t6t74D5oTk/w6uAUG/3XdlnC3MobDO5wXjWpWd3CUKL23mmQohZXfhsMJ4kG0RJP2B5j
ID2RwNTdQPuNVQl4EsfZA860xKJuFGM7kp0TOy9jxYYmDFCJo2laCfy9OgweGztgYkoylP70FMQD
/hEvb1ohEc0/xaqStcOw+FZYTDAu65YHygoT9nAzowFIIo0KBiLDJ01CxgLJo3XOTx3r5+AMA+PG
cNzX/D9GTmPZM3CdGPD/JDzSqQOFqvXEVI7BOukAaU0HgQe5quNEkr4Eao4GTqMoFpRPkoKBewuL
Qcb0NxM/yDYgCtC1FEqfsa/x1uSCYj5qcxsdhz+/drWOJE1/rKK2qkrCPOXg8XsOYYvtLGM/8rBN
wvPfBZuHryQSANUk+1XxK1xr26PEE7soLLd1rhb8riVG2OMPPjQndMl/m4muPaWwzBlmkpw0HtOI
l4mNuIIzQJ7SSRLes3TI+IyLtKcVYYItQ+bovpMQ37qlZ4J94qS/tyrV+k7+VyU/ELtkUX2MKhDZ
ayg1MK5w6FnHJr1RJGbHUj+/CSV2PH0enj+U0jUGxfQ2n/Fz88ofGvPNQPMA9gscULBUcr9G3/Cw
81gtiACYWCCp823VDBuKukAbgG2tNd8McCzBZ7Rues7z2PbmzjxKfKl7kbhOWND34t1G8M+e890I
JNCR6NI+NKkd1nG4HrlCA5BpitcjdHKq9R22Ngzxos4r395TKHpZTUwD12ViYP2iEiecFJfmQ0J4
nbKp5GdJpcT5riWqai0AbJ3O+sMgpzcFtxWFyuCk71jGCPLWTCa8OMUT1kY47xEMhYfLhl8U2f1U
sPWCUo3cCxqBcoH2/KMAbet9uFYLL2hdqR0bH3hAJ9L8qGMqTSnsS2ezlp9suerzIdkoymrODXrO
pJpWnJNZvFBJZmSbgkdTKxBU1syPAamspfpA4km90/T52vsjXDAYClv3pi9KxrZMhE3G3uSF3xLF
+Bo0ILK35b8CMm3OZG80qggy1oMOdzTozNBN6Te155RcGi3gTGgWdz5wE/kFXGYv726vNo+2JQDf
yvt6HVkMHTxSA6Ms9h7EANgnFaWi+GsTCV92Fnb4I4AN2DEYMCkY4EwY+IHi29cB6eYQpQglKx6F
+CHKJQMsO3Y2VP51d7nevGSp28zoY6obg1CqMDnP3Iw88HpqYtzJFn5NSLqQ26aRSe36eyCb/7R4
2yXQ+QOCUd+5p9FRUg9aBHt6Gg6zhmBNl5Si4DWxYBQYLAYbQZ7zpMXjOFYWORGantbNMmfDidha
m5ISLcKSA/sqA2iQw3tvWeFtSG8afyL9B86wV9SK55aAtwy2SDp4nF/dih6JTFFySBpnrfFDBCz6
0SnBxnlR70DdW5sXNpvRUrBhJ+N4fLIDp5J4ijKJCgelVC53iiPSlCfEQ6sCqlsxuQ6yoW1SyNAC
1JJv8bXzsqpnZCgC+6N7GahQBSyd+euICBYXtJGU0WpX645Cs8CrIrKt4M+SBo36BHr57o6gkYWO
FdzncGuaQKbVYJnBIhQknqTRExA+LkqyiI8OiLjeJVp3EFHoqEnfoNeo11HtPCUNB/n6dF8dVTec
NAyH4YPCACRdKJgNyFWDsJXHKa0mkEtFGV0+zNpGLA3MCSOQyLhxNg6749HR1Bm/xUBPVogOVN3K
ukFHva+n9gm1HNZjJO4ZheWsEOGRffh9ZIxjkjEcRo3ZrKdkq3LqnHka0Lss3yHQfxH9N2oWlozw
v1gVMSZTTkPLKEPlBJY7f0LyMikfn+vVQ7nS2kR2DLjAN17q5Fs+HkfFapbxIUDHDlML8iwootJu
100gj9E1NkSYXdv2xKjtXgSAZVujHIPMgsDreYrZNRdbhXb0PnOkQgqS37J+sL1y0/DLGbFxnwFr
yGRdPjnG/9yDNu42RjKwH6jsS6PWav6LHeV8pX0e0/e0kypf4YdEOT+COzVHg/tvvXBpR8ZU/wMS
p1sCv9BdwqZ9zWXltVfyxa7bmRiCQza30gMaQWoK8PmIn51t69a/JJc3Hh1yctQx4aUZ3/S1uEHc
MiYKe3mvmnP+K52vY71yonGcDKXdMHeEnz7/4OzzE/Tf7kHd1Fbv2nSOmFT8W4MSx6lORvebK13S
vDECShvMRCTvOtVDc7rdetCeCFVMX+7Fi1PZmu1y5UKbhUvkz1fJEZsmpWLV+3mAzCYBC+T1rSxJ
Se8ArhDBqbk9i16ZouYd+1U9oc4BAnG4A/Dq0azsFRf/9Fj3SnJoqKS+UzVDb0S7xGR2EVS+aqRe
g/LT5zu71qMvCdgR6w6z1beMkRMkCerTG+FEovfEM4+ppPFihAZ1WJxSqHRK8r+idl+NsLSZ0jYK
8VPo4yJbgK9nrBeGSz9Jre682onen7p7QNQxjFO64tg5W8P2ayeLjewVgQ6CMn5kS8xo3lawLEGf
aEjRhCdkgpNs/Xg4W/suacH+SXTGgR772oMzl3jxUkN+JFJrvjjalVm5nFMpZMilXYc4zpAr2IFJ
cOhUTcQc29VdclSqeBbykHHl7GsNyNRKAvQWyhmeFCq9Nfs/amn4dZiyHp9cXS1p1+TAGvT2N1oH
x0fmnD5XDQfydj+lb6PO+lS/Tad33l35GFi7oqL/qGAN5k5+B4sl+yNSMMf56PIQLNjylsXs1lJ1
ayr/MeDrr9pIqmgo1epzAuaCXhAzn/7I8+2uE9mN2VNdYcvrIIlQWe2cQsLUVzYEHb5pBEpPdFXR
UDg39Zsw0eZrc7bS7hQNRNSvqCY8EAtvaDrFzwcH9tVrbYYdGW3NfOco3SGn/kA7kSK0VUS7MQy9
aNkFKHA3TVleaea4Y+wcz1/2xXE0K8/i1Yx7o3CObrqJ4JGZtErBm+uJ32iG2oQ/2fxSbtE+XwEN
xBHWRSduULQAZ8jopNvtKqwV6WMuGfxKwDxSWD/lw9cfZoQ0tQQi+iPFPG8siZsQkwPpimXJP9aF
hNzx2Ji2dXlau/ga8TLnjptyXa8wyhk9SsV2D/NdEmrEgxyHfrrOhUrUaQExTM4TxmOH1oznRDVk
BOaBBO95MrTtM/lij9hs+E5lMs4BCsCufpNmND2ZybboAbVAYXG920/l2lUIn4TvEGHK/jEFJrIP
q4varu6maiZQqbiSxJjgyohTu4O4hdNjKVlmCU1yV1nO/H0iJlf+yVgvngvVf9eGPxxX3xgb7hjm
beIsXjgKi2x627doWSwbeJLm6migqbI5kUnbW13ZRrN/P4oEmuyv4PNaIdeOsM7IpS5h98bhNkNf
sEYtGoJINxgHdE/YzjFX6F0pj58zJoOyS0Kl712QLZtcpAmyBBAYKbTdf48gTdBE62/CYJYuT3B/
rbHBcY0OhPQ1vSwuCsP148PmbN6RNpu3iJPrQ7HXZKdMApqS1RGCi5nkNbVePO4Pw5Po9t7Strr+
dvkk/wmVOb5M3JHvP+JKTid6m7Z3UVC84+APH+zdhZzCT9n3XDbXkUvP++F1qQFrlNwQiLdrIDr+
3BAwtqqmxZKj2JQ3N/YpHBIlDhF4CaglwiBflSjZT6gWLnbZwYzTykF0JpEbrTmkzI/myh9P70q1
1ntWBZV+8W5X/cHAunGmhMbUChfkoPt/5Lz5uKOfUghcmBB8OYlobM/5mu1KkqCm+Cjh3++d4Bx2
fEouCcRvd6sJ7TsHJm/S1xQJtCpuzFmM3XWhxU5OzNxqYgYy8sRRVqLYBUdI8KfN8QL1ot/6kHAc
3TQWMcPYJ0k4wtKEm5pNtV2ixJBlke1zFr/glrdol//THOhwBaAdqd2mxzh6q5G5CWG7jxQ8vIgi
YzZCyFzNv4MTqJth9ORZxw0ujWllfo3NGbysOeF63CFSd4hA8twtOWEaypUCNbsT1nv1zQEdBnHk
MIBsqRQ7Zqb7xPiNcFu6KPaJ6I0Cuhpl3GWQyZrTSOrovgaFKDDiSdg2DCUhNpHkj97Ygd0MfXTC
Vh98O80caRsNjpY+Dvv2LNDQz1Bq1S/dnPoWnqxaH/oOliVtytDTKtk0Hy5CY+lSf13MWzm9kX/m
vOhjBmbFaim8kh10dTl2P07+H2dqTLEi3CJJ+RP5bd21xbtB7KUOjnTRvrIclJpdf8PLReSa7fFr
kqOfFf1G01QHlDUnfiPhzPYMFW5TADB+v1c3JqBG8+uQUlFtvVpK1ZkrUpawKZ7eJ3JuoUml9J+k
FDzd2tapbkkBK292RSHkTbDEbO1UahAtv4sYhgVy97HPskC38XC2P9+TS+nnKDrnR+rTcN20sJ5t
CgRh9LP8RaIUQTiiAgIR/73zi/nP0aijeXKDaGsZTq3q3wdXp42QHjxYAdBNqqcguik1JBlmVvbc
IKHUOGsaw4i0kNWZ+wCgyPAZZr7sxQycMruWa+FyOLZYoium8Q8AJ38W1xsp33VFIg4M/vBvadvH
kSj7zSaFypOZnm71Awjx8IXNc23l+epjOHOAC+MW6MvZum1CeGkVY+v4cGs58Wbq9/8bnBefgiad
vgnC6rkhyQw1VvMGwfNgGFg0hFirbxSt1CV4lAZBsuF3AvA5gHlYMOSfG0hRLrCHnWy5KKSgGxH/
w63u7I5JGn/yRt28baYhD8bzO8D36AojIl+E8isMgEFrj7VQ2e/xyFnBgAJLCLp6ZJPj24owrEwq
1NpQA2AN080V1EY10Dweks6JplhF6t6iFdFyEwJSxRkhUQyJABHyVbUAsb1GMctfR3LFIqH9g/2m
fNxYmL6zJwcAg71w9iPqWKAfb2nEd4mbH5OaGROYU7o9JtS5WqkwDVn7RBTley+7eeo5Tjy/FW/s
Y4DC9+svURhbuEUq0Lj6x5uutWjqJtPOpmMf51pogWp73APR66OjPnOeGzsm3KST2+HQ/XuldCYt
YdO1ta9gFVj9NiAosLF3+NTSaEPOEk9KIbIfHtaWxfdVNGfwcFfILF6hXCYT1WrjC4yoyMNHxB8A
nx2Y0786LO13nE/ty9iwKRSKiTm+I1ya+B2HtRQBBNAHgIV4xhJ7PTqU/yDFeuHoKl08owj7HNn+
CqXRY92uCOU+IcBOGHt6iM3aVHei1D6MrmOqQpLc/rTyoNkNDobws1t164EODBqhFABUUa1NhcgC
f2394f6x4d8XLN06AliBlpNezaWbVfISmhshT/ULgNwhdfE2ni7ne/SkFLimf0R5Na7eJ5kbRUMZ
IWpvESxXR69VTpR3cH0pmEIoTJvMx/7pXG72fEartmzYAcQ7UKjjAMjEi4uS96rxnFG+WW8CJXhV
V9FCAO9nL+BGkjKSaE8yCWzvN1osTpyNb6J4m9OtNi2+mpikz4iNbXmGvak8JFvd2q3HDRf96Huc
zO1Y6NUaul1VodaOW0AODN+QyqDBaJ+Gag3/kNtlSynK/sZeltikdf88NgubG2pPRS8j/SGWU1C2
WQQxSW+TJIRtbf7yTCwBDkdfekfNwCjYd0+j6TpRLjfrd06gLCrG66UL9jv2H6slKI7D0/wQvbvx
dr2r2bTdhI9qiBpkwfIBXiAFhssi4lEk5PcB90+wecVLTP4HydclCfOIQ+VU5/0WKKEQ7w3OgZtE
Dp/1S5TXU5Jr0pBvVZmGEBMx7J3piTTZoRk6lHapTxr+uzV5/zniXp8kMyK5uoI2RbQ1JUUCnENL
xYp82Yow56wEXHGadsmTuSBNGuYHKckr8q3zB+rZlk8DbIr8fgHCbL52VJ1Uhco3SVlT/e6M4wy9
Aa98mny4qTABapgeAG/VnDm0AENN2scL0a5hmwOp9QAS51RyByBgOe9VMOsr+feOW+WNd9jrSKc0
H4qrraO/t74XncpZ+A6fK2sfa+KmBqDRPbMOPv8BNOUlM7Q2UAcucQGsPBq2x/L/Ixz5t0EYREPL
TEkWyPvfCfsqudOeCR2Mj8ukmo7iWLnWZknrWbhmntBuei2cJpR9meqNMSCiY8Gfzekvq/l6G8tC
c5+I0A2uxGQy2V/u27Doo9cT+KCWhZMx4XltWXuOWJ6U3BaY3Nq5XiUnJpy4kOsLHlWQw8aGHSUy
j7JRG4wZ53pW8pfcShLeqvzF5CndiT9pxj6JGjHMfReRdKmxC+zzaQiSWAuAPc+o6DE0yFD4nCAD
XDsPky/o/lDg04gP9sPBDDd6PP7P8t333tLHQNJG3jKDXhS0Ts9J5QLCDJy8WcLZE9pjI5bB0n7g
rpvLlP3Tml1HQN5CYh9gZKd0hsDFYmGvsEQp4fnl0BNKXAELwZ1FQgd3fTJ4cX5iiHHLAOmODzzk
aFZm2zEQxnqfEauNf4uYFZcl7CvSGdpy/QyUQwMZsDVXsyQwRJtvPyDrzP9KyKX4vNhfir8StdI5
AiTPKMd38OAtu56tKNwjI9nFRdbTKiWy/gJoNA9Sx+oPnRkuij2KojkMNuGZjckB3Hf3IXzCPmSA
2KjsBBC5Luy3LNmcg06lr5rwVDcOtUMHrkpx22BOCduk/bnugRZ7/dqUOOE5pLILAjo8vKYDeJ+T
g5NxLuJYQNT2IoAcFDvLkL/HzFz13gpPgqLH2tY96Jr3djHjAGE83iW0CmD2/LhZpHOTn83fsdf3
Is/QlRuzLV3UWXizxv1bWBl3La7yXvZz10IbIAqG2YyfcHaxVecjadUngvqCXyyX+LIc74Qc7Qyv
qDTFeQfm7qD6MsCR8/tqmMUMSo4X6Bk1Xrkrz7ajygQPgxkN1OfW3x5yo0F1J+0DU2S4Cv+EBSDw
5R2omeX9dugMGysGcpXXi+WV2Kls9yYqkVFRkJW8HennNhFeOA7F200yguZuotlzrI3u9Z258w6i
WS2MXTdKhMgFc0zu8MpmysrtJQMVu3vdSZsyQhXo3CYIc7ZU3ao5IFZGX/8oHyPD/TFGGz7VF49O
2/s4WIKFijsrrbHNOMOXeZQIKRJWYSm0Q41qnTng3v3f1ceHRIqg8A8IzlGK4XolNkLueZKkRMlT
KKo8xQAvy89AwqU1T9o/0PERzA6wZzBkt0h/iTZJsjYYVGlZjZC1YLJ5aTos1IGMusYVfQXuVJZR
xL2kg+uekVk3Gn4cU1PimGKkDi7YPdFcpHiVVHlg1D7CZTJcklkg69nrL9grl6n307bYzcJYnOGu
NOUyoYNaw0kK1zfANLAhG/osqOyW8BL48KsCtCBgkJ8VY8b/lBfWSkJ1/HEFRZ7SfhxrtIyjauoh
bf+hawVG7JTOSE54OhpYswWCfg1iweqKURddA1Md2sm3qqTJRbWt01StJg6CJoP41mniHCN0jvTf
umeQz63yJEctiv+yWqOyvQqDZZ1amDlh+Wo53qYqQE0zl2NHP0RQFay/B/1ARHRhH8uQkYt2UF4f
RyqUv9426WJHrt0c6OMHiAfV54BuLx7JrZY9Zan/C+lPw7QcUTKTsZT9AvaRj/F1YLSPP8H9VrZk
ltNxlZa4FWj9HmJSPWal2frO2FMD0snXyfRkEhlpbNAp90j2XXO88T3/E3YYsZohuQKKD0hQ6v0C
YIg97k8KlpAmxuU6vU8FVUR6skpGnXU4dEB7WdzLXuB3szI2gWLW5uH31lp1zL+dzUK4749Q35NG
wWKOGNK3ex9KlDEC8toP47bAepEdHYycwo1NSvf5iylbDKEFvotxDF6PFGBszQTCZ2o4ZZQvb2IF
lq4j6iSRFYuNy+XrGRVJ1nDNLJW7dDSU09UTM9mWzFG+xar/IS8dK51P97HwwOBqpcoPjdxhbRJy
zJsPXDk54eU9xM5cNOEUL/VNAevfBNH0viy/VyluPYuRssiRXEDGi3QAfwAoGQHHQccmgbyb4UJO
gWg0iXeOe5wilSs74mdMcB1rtfy/FRtFJJKg7WapnCh9setg3VKHThL6qOu+wHGotL6WudU1gT7e
0cRNFIS9MMf4jhMQSOdnCGzILxHAxsO1arrxtYmOtHMkHjFBqssFr0eQrua87boodmwA56KbljVH
eoBjYDjW0ByCj2jO/YQmtEcQTh6piFLF3ANJUnS7i3llaABdTC8kO1zjZs6OIF+Bupsy6nTDOqqU
359jRfxW3xN2q5W8vK+SxTJfzuTuFaw/yWm8tiOfGz2BaLKhheNm/yro2FEwmEc9HjVkFzjOZoH1
Ze2voNuEgF1pd87EU/eev/EJ5vKJBxJ5fm6ofXdjAa5LuzjknPAJBqQujhfUNjiaupi491hH4Sf/
TBcKZLOaBqz6+85IHTHI3vexJ2yafgUBXlfYJR4M6/M8XXjEMFW7J52RtSLrIMexFBSVqO4FkAfW
dpUsFvP9zrOJQ+jhe8dH6xvFZ7kHq20Fdj0a7OGj4e7nJ35JNMD0smFlmnVWX/gg4PGmcvAKtxym
zNHt63GGhxPhD6qXeLJlWkWe1uSw3W6x/G+VUqaNcPBe2GW/nyBDhv9+FzeCzvv8TLgFzKO52XLf
/N2z4/7fFOr1F7ZBkqsBGhxYaeZUqn7WCT+H2kWLzfZD9OR68xFAbbZT1Oy/Vwt7/7Ce5ZYOAAvB
6cQygw4XxGsoUO9JqJ/zUfCCSLCnbE3m5XX/IenFWwOsdSa7n2slZuS01Lac5m4Zabpx4wERQkZa
I+7ttsBc3IuflO6gNgeBIPnZR62cq1bXr4p68MTQl/kLdUSHXaaxnL6ZGtgjqHHPwEZbBsGkJ5qt
lDkig6JEUy2j/xZ2y43RvX5KWrlN3z4wcMWbAqbtgBdiKK+/RzEMlCxyDSY/rDImeoI0PCLDk0Ma
spz0T5Mn0g374UOWMhgUnG0STvxJ7GKg52B2WLIMmUHtHEXXC8nUcS0Qc9oNQXyWlCEVkZIvE6vX
pnV2JNs9Ese4yW03Txl/vbSnQ7UJv42hdqosry+GUzP79cIw+ImFp/ma/M+W8iDRQj4v77U7yJ3O
mfjm5FY6Itou4b8RiwwZJ/HV198r9g4glIttV5xXn/BAugeAg60yL6lMXvAOfX+PyGsvX3aynEuX
pKDY0do7n77HW+3GNEaIcqKUX8B1X9DV9lFPNVBYyXLZqNyMiZJ3RZVuYR+NkQ1x6zg3yB9aPhDs
X6N8BXeUtTiWEFR8Ah9FTG7CUAjYluKWb7SfXWdQC8AkfDbQn97/jNjF93H6CC6yEZtcX9wyHxrO
WezakwoOb1yFOzMuoL/ok1YhH70sp/4dXiq2qEviWQd4jyjE7wcDCuDAjW6wRwE2eQ/Y3daRVosB
XAGU8q3qR8f1S8OMtJvcaKpsz/8p74Z2XNfdn/q8q8OwYMw58+oIAFVcDxUPGeNl+PI7PHR1nnjP
0iPUN3AhXEt9OhQ7AsVIgIdT366xbvdjEZPa4pSveaofwV5GtmMMti+sJuspdXCVFm3n52PZRDRW
kjWRi0t/tsr7RUOGCd+yBNiTiIIKKJCIOqzsYVZ0IgwRPXLyPwa5sn0f53/HeX0YIjKBtqa2dOz+
RC44iWC+mGZDGOv4uE1p0Hoyu8BTXHVMcUuZNY6zXJM/On8/iXlKW15UDXd6tZibP657gJn/OD8M
kgoXtMcTEEApoojW2+If0A4J5IsrIYxTtvhYh1l3djFSS+8opYuUVE56GkN/KjM3IUhR6dItlR02
qoJJe//w0u9e8QlkBraz6lVTKf+XkZGQuZF6hqnRTNgsDAX0MlZsWSo4xg5+JYLkHi2zZN6h+iPp
BtHB00poB5fuhY73Af6eZIglT9bhOROFBaXmKn0VNiqY6wMQcsjw7GXF6wRek4HvMxTwI5y0dVt1
abpA1yx/Shl9qli6DNZEYOYGEYXKhhLKWvtyH1wzgSHw7YRyPEgOAxErG0f8jv4OACdbfxxvTehm
AdOEMZzdUYGue6/NmEOWfJQAk6kT2pLfmXGMebRe0xSafU5RjotIqurjMFmJVTlBUG1Nwegr6VRv
d2q+wy3w5Z/s26M5/APlHnjNJg3uDBnCD7neorlAohOBGvu1Gsm2AcPYhiRK0rouh/QCVvRcHvql
3x2ns0+kERRiXjh20uVlNtuPVn3ZmypS7JxZX2Lf6bcNBZQrDtsMifvZJos4/Be6votQNMDJTjED
924mCReM+6R3HE4veTQGPwJf+dyWkpkrcMlArsIJclCXLhH6LPQvQo5u51ErUVdMliKmcZVfs4NZ
mbxBsj6FUMoCjYuLIBty0p6A/kt3PfqVuoGz9SLC8sf8TUZrGcZyjUcfyyj2NoMiTcXEmD9gjJMg
dBCSr+Z+EqFNcF7Vyh3ISieb1XKqlQim5+kH0wyS0azrPjAs3fA8Bw7q0d/3m3bpOhAQ/HhdBSSE
bYSbEcfNElaUxR0EdoNrUYUymoV1Z1NI/JIXddtayp7otNltb4g8Tg+1XobTtHJfLTcZpgDXth3b
/OMw+Yy1jEXlguFJALtROewdJCN1X4akXaaxLzkIvxmTU/7FsKDnuxlpPgRESsF14K7dLkcmzTsI
qgf9+vyDjKe0Avokn1G8b+ZBXPhm8KbehMWQOYlemiKTSCCNqTkurtxAOfJkdEhNlnMcD9ac4KiK
ejm008vgeFDft2avLvTsXoKGwTerCIjOTzhjQhnSND+Gwjf14hbgvImAU1jSVmPreW3XUgJpPjaF
0+grFseVrQjyEKNwHofa/4M/vD3LHI3Blhg6Cq4JFoU7IBb2xIIhwzggZlPPZUBockTPlIBpoZMv
N8kyqqvfXVXfKwtDFtdUOl2+LuMZcQdhtLGsPe+b/pGuiSej+PS9x8I3nZYec0mGsqLu4bzifOWV
K3AkPCh9PkvHniYdlc+q34mlJRQn44yBoz85xV6E2eEj5FWb7rcAYSEC8nwAzRbCzt9oPLZRWGyd
okTRBVys/qDdZvysVqHLztxdE86UkUpxPgtdTxroe8OOakyut5s7GZSAW2YwY8z6ilYYp070NiSD
5MdfRNRkBbJOq0X2cQ+T9y/UnDnbeAHBdlVa2lD4BloeUIfUYQfAxNmghWV3h/VAV8ieW1xCghn0
5apq65RCYwECvU7pVlCuKcB89/s0vFup8FTr748oxt9RceZm22HeGr8llui7nNdZw/YyPx6a9ujk
TtPXVqW2GotwD43LLC+oW0OuS5ShIUMtdJCDIAN2TDYO/Jm/V7tyNmRLwPARWXd8pNRJmHAXWM9n
hHjRgVqnNg5wVxxjCk6nGymZIlNK1Y+lZk8SORx+xWLGL83dbNvYSD4UdjEfMwekOQPA3b8f4dWD
O9lsgU9rcCo/XLo35/eYvNyrwUG+uSXvPivoO0V+Td3PzQn9IJ2X8MhUGGWvvdDEStyRT7Jmupjb
L5d1UuHHUwqd5+VuOHtW8ad8lk0dzpaHiDPpy4whW6QYfmrpnsaHufh3D6ggvWIj0q1Oym1IqhOr
sDRQ+ws9dBNPG5z8fGpNAmBsK3klqOkKvCZRA6mz3re9NgDEF0U8ul7L5ePO+X/CIg2iFuzriYOZ
TeaHwJKBt6Cq6qq0SEwQ8JJFNmAE7CENHr5OruEcK1+ibGvWgCN1FLxRJM490sX7okDq2B8ngrOI
ykGkf6mk6dH9UsnzfypaupI8gxjfqYUWf3RpApBUTErB5yBwSRDPVjg7L+tTeHyLZl37WKhiDj31
DxbhtX97pA8GeIK+dS9hbhMUSCwFUQPingURnedYY5B75O8W+9HB55cP2hbNKRCh99il5ys2TarF
SLOMOyXgN6+dDg3B1YC+wVSnsGUcn+Ry2u35/ZWppqRnD3u3ToYASU7p6csSVEcecFSbAfe7TK4s
0Pe07lAT4NjoJHfl4vi56liIkQY3A0MhdUYqW6ixsytszqqNAsnAch95XBN2jmZUBea8PMSbK/Iu
B3p2k7WM/hcLBUs87z4IKgcjpmtZJzJUbkTFJpXC+f0Vpv5d+5jIO3sSFtF2z7nOXVEoAwmhCPEA
prmDwmFFOEfGYf5EuKVABBEO52aCUhsGwrm6iD1hAmLhW8ya4khS9udhJCecjkIKPmcsADSNW7ma
mantaLA57yV2ARWBYQ63Jaeb49QbyP97ySBu432OF6Ozdb5kQiZN8NQEuPj9CKB8nrZoHRHKWjRC
B7ui5NDUmu5fmCd5bh15SzCPZxfxf2JsqbCTVedJjhA3FqLzCgYw2tVZAgag88eWmLbeXQD/o692
B70bBPqGihGg25Cm2PKspeYZpIZWdmeH33eYCL7uhWAL6o05gqp83Zw5+LpKxZ6SXaxw3GETwWUo
bpSO73K+lBgFe2nNV9FS75I0gRO8FNEFbB65Xhq8Wj6NWuMS4F4ZChwqsOUYkh5/s6hdBFCb/3Af
AUeGW0mgJXE6Nw821rBIhwprbhNPc1e5DKLwEwCizN07ysBu1ej2l7eH5z2Gb4pgqMrdhfdYI7M6
/7EoJHBS34ipQ4YYx00hhQmwvGA6tU0tpzqvSfcLC4iMR9zY3v2rFEzHwq4uVqU3tqTRljK1Hs/g
Q1tc68hQu6bFxldfDB8wZnn6hZBxvuJLxfP3q+flYrh4a1oQeSFWrkt+b+24/V8oL/gElDTxn1QK
iLRGZDC9cthKx6+bHM1CelDUEJGv8znj/Zr1pl+7zpRGtL9MaWsEMgjj4vhYSUqcUrWZQz7s3Xo6
f6ech1d7TwTVr5kU7C6qAZbU0tZH6emiLWuoTvj14yVnadnYpsNnBgqEbsiJVelNgaMHE3y9jKRC
6NB2v/1bRP9RA/A/SPtaiSJgw4H3hZCwnC/1wQn00K4NGkGIEm465DD1Q4zTUTpnCECfyQwpqvYO
nttkLlYUbAyzER97SJL4UzoOA95OnfG/fag7ZQVqtXIBCMQJaxew7Hflb+S7LRW0VdxDEkj4lfpl
OcF6FAXKuxH+OsKeQslhfZ2V29X3PPHNAdmzop2ytR3++v9Crp+PyT0CWeL+lNor2h7NCA9dR+iv
q8VDO1bFvD69Vbtt6Rt3ilT6tRIvPNbWdSwhN64gs2uiQLELhLPTn3XnTU/hQ+NFAufXN5F/bEVe
zP6gWPif5Z8H05YsakPcAh4MGU0xvfpQEUkfWQQKM71t66Ao1+Q4u/9LFRQ5I4hZDdetgys7wQMt
3kn5Y6h/D4I+6xy52bL1vmsW+/OuNJTwjDHHMRh3ulzUL093blWkE+TrxPW6k7t13uaPUl3QR4nr
brJLKxN6ZarhYzeI6qDcpON0JIgL0Pr7IfjPyI09PVWpzehnyjlLK278gnkQy93nb/xmkOiBrKah
JgPrT4nWw/4r5OrfKu7UoiPidC3uF+WSZmdJcQ4baijypahadYLHNY10ho4SQYD6MxNgda6c4AGD
v680Ro4NKBm+xYs2O86KD9jjIeNjDzhN7iprgjtSy/YqSjy+XSRbUx3kK8CC8Vu4Yn8ucI4cRqkC
N0tKtDGxv3sHzc0pzS9g1QY4+QTYLQwOoIoC9FIkmRuDiMIMiwQTFqYHvt4z67bLe16vTj+J+uFo
IcCu8w96/7iAs6Vvie0obUaXnolbFA1ouXGQRXFq5P4QKeps5wUgw0YHNdNaLGoWtLFS4oPMZpld
Xlk/wt1fXDZIdVEEiuBc8kaBIT5U33SMpRQc1SS5aAEr4YtVeDjbOg9+wi1l0CtPgrNoOFrBNFDG
2o+WiIYAGyFny8GbIi1hOqpwY4CfbaKpIqMykM1iRibGFWd45tTvIizZouptIDQP0XaIPEvKkQE+
ZlIwU/PrMYHJD5E5opKa7ud6uUdf1wmnhf68NYTqYKrJuva5M85U4BG7Ba5S31MGDosjbkY2Brh0
8kZzRdP/dzOVtFTVW4W5dE0tbmlJR8AHbnHXnz0YE23b3jPLc3NNr5kkplgInDSSNi+kreiDR7ju
vvEimHRyykeMakfdaUyn6q5Xmne3h64wAoNY+JnwYakawwCo44qepKSvq3ou7YhijHQMLfLYsxdv
IvySvH+nkllUwHxtQHWGS+juNNIEEa2A0uDaPIMQSLf2J7IRa4nlkuydDJNBX0RgdVgZwNjTRmEI
no7nBuV0+qhlztojqJiqT7SbC/28DJEcBxMO+MDESxh1iNYqLxzsDJ2Q6hQA9u7apSsXDoSCJSpe
VhUNsKkwdyZe9Q1ik9ISSbHlo3kincrR6KLUeztCVFG9k5JyKKEpKgxFP7aASGiEgf6BU2NXO/n0
QTSIHfn/oUTwiVDxH6aAB0BwQNGI4QrhlD6dBL9Li1Euti/8Im1egbV3IAGOHdJYyDiLkyDAC4Qn
TX0GhjXsTDslLX/FfaQYKqrLoyc4mwHMB7VOe9iS+27VWCVklk6MTX9IpxOeg0s2lkCCRkVkkzXt
ltSI7mCiZmQzVMQk0QYhkSOwunhmdlzHbwhRzYOStLlmD+vFhC+qC8kbEXnOcJ3uLOENznzOTGSN
ht4sB1n9Lug4Ripf6LZFDuFWn8SgluNM0voOZ5eJE+1GxUMPaXBIz9ZkQxFeJYF+tKmz67iE7Rlb
rMkGCQzmIL/kvpMI9IyrE4lZK4Nof1apEAqhB3ehYAidtAgmwHkS158fMobz3MZe3eQvkqxu8XoE
nxC9xw6xcsOeiPbDEBfKbzGjGtBNns2hc7ZIwVasC0LmSEvUvtxMRF8MFr+LE8e/6fbR6Xl45rGM
MQ44XerKXhEW941WOBfsDKfN3kWMcPM42M5dCBjL+MdfwjIWA7NsRPyq/DOqvM3UzvLzC3f6iwTg
7KIMUqDrVoAaYg0xiKb1PjGUNouw0bZ/Bhg8zx6WJi6KlHmdL1OPqWd4QQa2l2xk/JNA/PIUL9w8
wj43ZQdXlXccVRzMKFVFk9S9p0rLbahTHdnDOa74ay5Hh3ZJoQ7ELONCSRFnkszUJc3GTsmCqK6b
quebjtovI1p8YXZJLPtR1MPImETM7h+C4TAyT4WQXxuK1KFMVjh+LbThFxTdQB5ylEh8kDQdnkYY
p89l7uOpDvhIQcBhhwdBswj7HdIBp8mqIGnuXPlEt/LMxbwtyt+0lNDJ8xrkFXpDUcqq/TiIeHWK
Bfw+do4pD/0H08RQmvf+GemGYGtktUHhPobHCzTBHuEqDNVItc+6lfuIWe55vavfCASnZ/H6IEGw
FCO2f+j7uIuFgxlTm7r2bzOQYnLcXEjaF44XUfbGhOF6YfuN291yYc0+HWZEHzhzLnVVjM+b+okS
+oFaGaUhcbh0L/+qpmQw8MWGPDrxP9rGjc3/DduqhoHhoQXtuo6VtL4PtyuEYW90VaPCz84NMzTj
YbMdj9SR619gagtUaJeKZUneW1YFWjmEjMopHdNIgOMcDrihMx15Ub+GmajG/1Tjz114lsZ2VXjV
bOVYnUao92bUGdFEvNG4ZUn9Ik4bd0W+5Y9C0IzkgtU1U0qh/x2R/eQhSJOqxj0iLw9bnqKBRGQ8
hV9eWjPWytrO/YsrQqIK+lk6NlNs4CvKtSeuTm2Zw6VMh4MiRSO06zS/tmmUp7uRVtXlvvw2oMNE
sM/MzkBDrB5vWpuTn2kW0PetPT10qES+mNEX/uYibqWlZVcdLEIcd6CmW1LgSCDHJ4K+UTeW4k2C
EZDXunTmOX9TmGuM2FQYDRnN0b32im2IeOImJlaTmAh5Pt6Q/A/luqSrIKbA6wfW0+8HUtYkmJOR
Qr5xBjcqjVNZIESCqxKu8vlcWuFZzDMp5z7H4jYfl83s/514D4CkhpaP8SehOf8dp1B+zrv0OQBs
Vd7ZYMSu3rDHx/+/WSBMSf/5oWSPZRzKDQZ3EfgGdEJUpnxi+CxNvmZQOXQd/jOgGjWVhyp4dkyV
aOwQe66ZzLoIxijBLiBlcCekLt5lifPFtbpsuS/gYIUlcrTbyDTedulIG+P2qswou05scLAPu2bw
H1r9VzHob5k2+Ag87WFurHYGImUPpTpmnS6FwktXdO1zToW+wVyPt4wX9MrHy79vBgI8wdvCLfxt
eqjY1m9ChgM9pfO+6xKHVcxAsRLAiwNY7dWrK/eHDCzfNZtr4zjUd0dTfXDMaG0JjvmmW+3V6FXO
s5M2q1w98Oki2ZCJtJUfLhq07SEVhDUohODExgfeqZCjbHWYkpYs3yJ0dQxH1uZMPgkMGV6hMFdV
B1ai1HvGsLntwxDzzRPodYKIwkR2rLCHf1wfyPsnQ5qfAcBBhrXDOzKqXk15Jd5rrmfxnoeITZ1d
mVW+EHa3nMN8Jb4BcJt96upgQvKbVjSLA+sy56v/qJJiukE5gqGLqLuDCk1fKhVYL7cPKNZOh21W
qF2rbw7WjL83YU6ADPZtaBKzl3nJoD9i+BJUlES+8xdeDgUbMVziZEH5+Anp309lt1M+JYcmpfSm
gzDD7VE5k3darVqzDPjTgd+6MEIdlNhQ8gaM++fg84hNjjAV7Ea5ko+y+cszNOwNBbWw0RG0c7tP
0QfLsym2WdjV9M5ATP0pEKopv64CeyC6A7+0T4BjTFo80I5YpwNSY0wxFz2Q7fTjU6WJ2perP0yw
OkdLXy1xcYaT9A5VPUwhdiPE7dld+21joO+y+cFvldEGdBAeIGjIe5y/+HYdCJZnJh7O8Z6ZNl5B
LZ2bfrVt3M3v7FSaxaxWKuONMjRWWyZC07uBhwNOno8eiwnKElhM301NuvRSiBWeGZWjRdfCuM/H
f7H1gzd3zsqESZQKYMj+nh55+mByE6u2iRIjpKsnvoh5W2OhMihIKShE2PEi/qzJnCFFss/ZVnWa
P5MwwmZ8nTFEev73K/w6zZ3J7g/6RdmmwDZuBN3dH2DSPNtN8HoMtI6QCfE93dLPDYQNJZysR7xm
NVrjJ5pu+8yVQwjqadtjSaIceaGz50peCSIRmBlKSDFvJAEBB0gQw6XU1UNtySvPgIKxaWtuSoYM
q+OG+NyKdpEzb2k9As2HYPeHbW0279Z3rSBxioIahuz8WAJvL0N0gopknHiTAuZtaKxB7virU+nK
hhKhozWp7ZA586RmzOqeias5orHJc1qFPJNZuV8QyJ1hC9dKtuPCCvA4S4FMUM2Z8Jm4kDOmI07M
LhaHxBIoULIs5ANofQa8MwuntMgMaxfuQ5H80Xn5wwV9Dge2mGYR0e1k3Oa8Ul9h1T6IIlBuNG8r
5DWYagrwfUZipqmDI2zfdF3pbqsHv9uku5+iBM9dEU96Vws/8PdFGfNAMKUfZJ8UrCfIrRfSA9s0
ZVV+OjQrjS74REs8Io+GaUMGmZ4vTQhwm0tBYxtHLCwx2v4ZCIyvTazlKnreb852VGyW5CNHnQ0Y
sohHb/ucpOkFnNTgPLkB+R3iT11J1/B+HZpDx5upk8tel4WkC6PzJ0gSdG7GaSLVG1BinoOXNT/P
iTE1WEqOKrIsvRdrteZhEhpNY4nfAVlIQdlhfIcDX+Rkj2vhnHzxnm+4Wwsd5GTfKk0dplYBif4p
Igj161YaUYvI+gLC7ZW76L+u58/1Tf81okFTnTRoiNVAPpE6Z/brT2CpGOIPo0JTJr9DpYL2ddlW
btF7tjQ0Z6Ne19nCxCVQw7GSSzeZ+mAabN1FPrX+7GO5kNtpNYZ8A0sA7vbc3HjPIbb5nub2QGeL
Is4fpEi9vcgNf1f1SqcEEgfZ9/ZwmtN6Wja+Piy5f6oNjgfIFurdKIlisYhiOXXFjIjWDCFr1Hvf
5mfmnWGfRRUtbC3e18UAwP6tJBOQ9fMPgVLHmg144U4Rl+UYDcGuuyYxxP05l7KtCpVoqY53oKLM
IisSmYZEPplrwnF1hmuRUkl2/D5kGZVyv6+sJF7qnbr1uJUG2rJf2BU3YSPy7+EXtjtTc01t5GjN
kLZXCkIYIYbVTe5Uzpn42Cun0bW5EIb1cgzX0YB53A3/KqpyY42ECj2KSJJgBHIQ7oDY+vDI++gN
FFstA87reBAQOLlhpSOgDOHemWMtalWW84fg/unOnGq+ccE52aVh4T0Njn3oLHD/G0QLJTP7XNL3
Dzqg5A1Rgpn8dJTu7SUitINiua0I39LH7N/BZFlPA8oHgf0jjiKt7jnzKGHMaOKSyQQ+q9lSOTDr
2rJusOWuwNf81D163pxGNuY3bTix5Y2PSzvjyod3FEdO4e6tQoKAdCJ9U7HGfkC5f5QSXRW66cHl
MOpVq7ywZ44Nee6A6Lr0GSrEoAIHkdstdSHcEO8a4SlmaUcofbV/UHMdUvMaB8b9j+WGdl9xFoYb
ah9Xb/yqOLcLiNyovYkThwUT6gl0OYhcRIcausx3V5itnZGh1VvUHuTL1I1i1XGneIOKPCT6b/vr
bYbiFql7LzvGwLBT3+x9F7uMMdUTXvwAIrVgeCScScLq9eNroh4Tecd3dmYiWMGmEoGKLY6ygE7/
MXdgSkW9qxWBtZe6F7d3atOdauHy8ak7VxPluHr1KI93JMd+aI/uAh0IILI/6EM8y6RWH9y+k3Kw
ahHEM5zAMq4hmOlECIbQdXC0VGKikuHhcNjsdi5tEgA7pqL3MQjTyt95OZE7DUM0SeEShcSYe23E
Z+92UJh86F3mTaBnyKSneTOxuPPSuwEq3hHtYTNARymBSuU26Ie9+XCvb3SqSWtWTm43uwU0WJ5n
xJOs2zTjYKLenhuUFWmIGpThlEzHJw8/Rrmaq/D9VTfwHjEELWZeqpF8qwJfweJNB5DjhdNG8AQW
rxkjXU2HmZhGofjFOKxbQ4E+UUoI1/HkLtCSRXcl3YNdFdZ/r3qxc8HPK+8O9mxyDCwghKG+rkuM
Uh1y68ftJITei4cI8lVcffqMPwf3qQ2nUJIsxCAuFJQUSz1RNUZU+sEf7mupVgpquwaXyoqhERju
TcvlbvRl4Zv53EZzAJbeLS5LfSH/bPmN+TqbFKR0pGhS9a954Hlj3goIxUBEkGrI1eiFg7Li5NVh
m4EU2FvYVrcxkbEpWpcxVQCDFVTj2tjodJ6mh9n/uXADN+9SxOeeLHEkD+ZutAIjxOij1+/BLJUy
5AQMmMXxpW7nZGb44dJDhngYwbVOo3i4T5T2jKIoiM6rKj0bbFEk5XFs62oD2ZMuMSLgZSoqMAyV
vrqtXhSGCFZ//KXeZbawjh83HxJHYJdRC7L1E9GEAyIabXrUrBeDnQLQnIGU2GpuaRmsPHznaDh/
Luc6LaAvM3oE0XHaKdRtWWgb3I9cR6EiG264sL09pJwv5CEWck+W3WTE5//hD3CNPWrt0cYKiGRU
+mwUn7O1085FNk/0FPdKKajqNaAtXYtx4q0WYRAg1uetIZGXlIxvA4ioTB9gt2HoHYtDh0NzVujE
cBqPkHPwu61uuy1woPfzqIPJhLki8WFg2fP9+4XDp+1J3tIPsExrAVsslQ4S2cPevJ28gZnvf8he
c14VZRGsTnlUVkzvJNn0dZdZ9aJBQdChoIB9C+Tdhoczs/C8aALDAuHS+PBIPhc4NlzkZWAo62Fq
JL1kbvFtsztni3xFNhaUq6CLyfzSdJ+5S2RGiD1Qm9aM3sRZfTa3HazUMlxFsfVIY6vVf/Awwcjq
r29zmi1dHlju9LzPAMxA+JSrAzylutlS6Z9OuvWMKBURjm3N8pPWBOG5B1PjlcMEVGhKpybb6aUM
6Agtk9SwXyQCFpE2TCExOm8KZAaVK+ap+W8OUJgRunamTdAAjsGaC/18KaBd19uP+J4AnFEwmIYe
SIbgHLxQNpJet7j9cudfI7NC3JM8sQerNPz+zsSbIJu5h1ubLquyf5snmXRAki3DDQmWdKDYNGqf
pM4Skxdtbr7LzpXOpecipw5SecSOEXO39jHrwvgWJVwbXYE3r8Fl19k1Iude06wkNNWTfwVWz9Cc
LSSXoN25i9rp/J0HN7mQDT39TwshHGgK2lk1Gas0q9S1l48Qw2dcNHOEPeUShGNcxtzIhgiRJe6L
EyyzYIey7jjM2dc6i6qkJ2LB2kLJXmvfJ3Ltb75ad3PdRhq8HT/2zHlCxazQ9BBskLLzj2AufaJO
Jx7f2wnkxXAO6pWFchzSaK4RrETBAM8lV4VbzYPRDuOT9wvb7WsV6LpUd1gtniECqnO0nNVR/5B6
8Eprri79DhkDDkyBbshTXFdBrv6y+8Q0ImqNOTQYyLeQd0S4ZynzqCacVPzeI4xPSnHdPoGPY7+S
xfnJFbtVV2E1TsVjsrraIjIpf6ss/FX8hpRmdN84Pzjn/QID/IeT5kR2zcUC7tX/WmYlCK7ailbf
qf3RXEQlw9FYQ1EtT2qENPLb4/9jU8TbjbEnyPClyMwfB2fmFBWRo+zCaJo0L0W4ecrASr4cQj5h
rKZeuG35Aqrl4pshrKAWsOXIgpcJvkBgPhMRq9LzAITXbgvNQhWpcGUZlgvVLqLoDS45B8zvxjiN
/uEZryH6sZKVhUcr/9gC5JRuKQmquEm44zIrxnGnuBiIO196DI0tEufvCfB9vj1KzqKFn3/z8OTb
8Vcb4i1gIJbRBMyNhyLFdbtpFFaJwqroyEjdHoS959qD6n5NJIhD++jUdoCuNcnlMLdZLK9ZB6zD
KOW3fw8ETYtOMcVZQOeE5plys67kW6tQjQNU7auekG1ii0ucrrTFTRTQWolX88VroFznEh6YRIYd
v8owRMIPtHMtXR2AmeULNGHzS6RvX3DVOJE9OOUJ9JgPwNLr0gU4dY9ruSIkzs/IfMnvtkt+4Bvk
s8lBMFVZ9cCMkH+tmNKWTvJatO9yi3FbKSKTexK+XCqO8/UsG86za7ZasGvQxfa8rTscuJGKHJtO
KMUkojdNaIqVoms9eRdTL+YofRou7WrpaOi1hPYL376KWYaTI84cZFf5EGF7rg7Uq1Ih4dDO8OLo
pWH3Lx9my9HhlCESIHcDCy9yyZFcW5hDRZRP1eZQd83+mVYJqm2nkIEuPRMuA0c3JuhumvlSeIP+
pW8eHOurbZZ4dn+V5Tl/MPG048e8kTvlVS7TA1bzyOaiV+QplvtO/LWUrPH+XMSzoqaHcU8m+nps
EDY5OFWmJjMVThjgNqtORXRon7xZosJ1VNA979dtY+v9oM0RjlVtz/Ho8Jc50mEDAcWGBoJLSCdU
Yotybc+T5mxIglfJnJB3jzuHOCDCzdxjW0XVKvCEwpdiTWchw6RcVTbfYE0RkPtqi+RUrLlluTKA
eu5xnZ7+XiX5GpxuQ1G8k2bqThyYFCNDfnrJXg1pkKcyamCdNbIOc3AJ/5QdP4wV691PRTVKilds
QbGRbQ2YZPHyqaP7IoAr52YQwYCzJWe5RzQOf9O9gnUet2yMUXAiX9ybw2SBHxB5NzSVFG2KZTTQ
rzJEfaEYu1XUWJUzCrXX9eGL5UNegDI9lXSDL5OY7q7wZPoqcCtEWEsk/ZGD2eG/aP0y7wn/osbx
opfVNkU78rBkn+Xm86/lZK3MlbzslY7bWrJvZtKFxQaqEJ9zizpF4r1rkbUt7Fa1TqJ0eBeMpaOp
NeZXEflnAMlRXb7TRNeTZvuUWefX0cAlLJKmR/zyK3XAfQQ+gy/3/+fCAFYN+sjrBBJ0m8iDFnrb
sRCKJ+4gvvW/+Z+tkv52gPpYHRtUE3jRKvbCVP88e0deUl6BYj8GGXMzbmoOGhAU11LLhUi7onSz
E8mbs7puGagPY3LTRW7Ql8vDAL29FrmPSrttorRhcjquDKLL+dkoD/ARiTAeQRvL1tagy+z0ukMJ
KttaRlpTka7ikVcQJu4Ovrq1MuWriz4h4cRCRgCT0gSFaPx+ymKvTe5s5mKPHKx+lOhChLQow04V
4Z1WAJjp42guBn/bNRBFVCLMkztTnshPF+nK/oxg0zPyDUyT3vlChaXoy9zkKJHgXDB6aXoVNMCM
Tty34hTUpUubyFgWZmW8uGfrD1OCL1YtqWNSuU9INuhg+NThBuoa1Q71uimV7g+B7cgnP8TcKaQU
OS74hf/obCcazGdksKnoHGnyqmZx2Pk5V/DrZayyLC1n09A8L+4Yfl53T9Blxt1gJ2OqH6d5GWrd
Vw93Lhgzc784/1lmgUFJClQKU3XVeWyhEJOE4DKFlGoULrmaNmwNeqdMJbX4EN9u6px06EPQl1V9
oSwmS0I36u7DP7c1lhMvacOXU+9xj+qIYarNeDZZcBW+OJJ09gaXyv0eNvuNPFBRSKvpqJFR00w7
Here3TKxexkkdlBubZgz3gkDY+5K6+ccVov5qTu41AJnkxswMCXOVcQtdNZDx99OQgv+NSSh3rYM
oRTDSTIqnTvgGjqD+r7MJT27o2F9m2bufS7LTsxPsQN2V5IYEtd/Ix5wZUPF3euzLT4WMCSkFADZ
clh+Yj8/goJD5e+y5H+zlo744CiFCVfh+milN7qNy2xl8QJiu6V6JIO7nIo4J3tBKg3z6SioshjT
73N7cVrhra2hkXE/EDCIKGASzJKBuSnBWiw9TxHcLpS5TjiRnFW6tFMXaI2SWu/tdRPZNvS6QaXD
PKGyvqi2vP5biYHXd43ljlBS1D2KNwrGXvPp4pMZKwBtkeRapF/UxKzvn+sOc6yr7lA8fcPflqzI
USV4DtVBFV2o3y+29d96mMFFtYUWS3oXCuHySxADTlBCNbdrUxFpmlJidcEBAG53VG+ldTrcJn8Q
NFhh6kzOJqQZoNoRJIW1LKmpB9Xyn8UuJ5bPW0RyAPsONc/U6YmHkP1Mvm7WmcZPYOhxslRpr2uX
qvcOxWPaJ+2M1/bP82QiyL7hihp8FIx1GKMWnUILbCoRZmXVzevgCZWG0nZD6dLhPek5NtmCf131
aabU5v9zlXFeHzHDBKSZY/urNl7hs/TnvUeMaQK9lJI0dqRHUomBSSFYDn2VNQElpZLCUh7Db7AR
BEOmLhxnFMt273whjrzG+r4n4pSt0Ti+Kb7V57cS9M8U2WlHvcwT1LWktQWdOHQvLL7XoB/sOodt
9n181e9EBL+9Y8LbI9Ml6rEybty9w1qhzMJn1q5zdy9yO6nfsfyRkYIOyzUDmg8OJ9StNuaLyDyA
+Cf+mBVvXBQQz9+VW3Mh8QTxNqsTWmg/GbRCYWyuem5EybL+sAQe3HxtVjsFC/knupIU8IKJqwVq
BDX/xEbkulQxLUAv5biSPZ/8UmWWm3pewPSM5VUQnZi4T6jPJTOBn5gTGJ/cHU0MzwVXCxvatisl
oqUIOBaPrEM0j5Ce8gfBsZNd0QIj2fen50ICvR6Xci4LPtGjd14dFat/GSGhRoHk1B6StLYAunvH
nuOzIJgrmlUfvYtJpDFPBrKfMshtfAe2Nt25dHrnaD9GWsY6kc98Re9mesoMPFMq1IqWn9NOBOaX
77BGmVhAnwUsjq2yNW0UGKtD7a71C7G/9rZWyqhHWpm8qlOt90A3MR7We5VHUTqy3ULwWnc8XtBU
1p8PsOH7q87i1O1OxVWL6haUJLY3M0Q8yWTbmWFddom4XojI0om4MFHtUiDGVFdOb85hG29YcCCm
DU8OSWk0zZqYBgt1MQzGc8yAcp0pFesulBeIF2dFUc1HNrjmu7usDpgArZYzuFl2mefDTC2ybdZ7
vDAosq6vhywWTuK+hpeaqN8ZXpMBCBAqD+/aaScoV/qSwlSrvE6O0LwG4IrVX+ipgNjG070Uh0BT
arf7oaELcbyGCaD1gbbYhqHX01V7ZVX5GckPZHzB6b/qkx0IJgqFjBxIKEIOGr4pzgec+i84/2oH
hICuTJqTa+qM5FlDcf0BCcXIqmkG11VmiW3Qf1NqHa8Ec4j5wCyFJbD89BZvVWFXD7ByR5IgSS/n
1zhtdntIH4PhbYZ+dXMSFotbf5TygWJuMXJgjULZ5A//ZAK8uwbnIhHGz7vMoR903bezrvUnSNTl
JAGrOYGKWr40ESMGvINgaffLLkWJVXnveTUl9pHiSz9t+RRR7BJpjR/5WsLtg8/Rz32pW8T26w1A
fYVqzrkZt2gDU1TllcmRs88DYUmKfiggjIp2d1q8sAnRAnYB8neimffNj9kmRas2lW93n3IzH/S/
GsoKNlvz4A9oE2XPG6W6H8IPVHKYaQEo+JA0MuTrJvjV5cjhpRfyYmMhz4aKvehU8tklgtpih38V
ULZsEWm3dfxtfliSIGbvVGa5euNLtDedEeiUNgNZ7TgZGJjWKoRZwvWP+1miRpisUDx1V3gTba+N
zID3XFo=
`protect end_protected
