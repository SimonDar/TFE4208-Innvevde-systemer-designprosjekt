-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YndCA+B+LHLCxveMdqwuZlU1KAgeIAmcPTNQVZhfzDM8ORFor1rbWUUpS1FAMcWZyQ64DazyiCGP
MzYf1Etz4g6Euods3OFRMipHDLIcckuIo1ZhFZwv1v8gaRWDWmTHEQCYqPrRHTlsB1jveXMf8j57
7GPI7pxMrlqhPFnvhK1v4K6MiRlcs30LPqjdnolLWF6ZWva6pGhkgJrbThTT2glxOu71oB4+hWRH
jB0HtWArv00weU6t5gefy7uCXUpgmMgtoiHJB8RNtY7qGFuwTcac8vkpTnBydBj6efEVR0hCW7wQ
gPGcXztWYuc+H+4DfByxNGkQKV+s59Z30S1Q/w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
rx7vNywZd0bZFtjOCXGTSgJ9Cq9TPmfi0w64M0q9g/U2F9UQGc5fBbBSfr/kHQHbekmUmPNvqa7W
7J4mHX3f+NAvxkfiqjxGGHvunOZGLZQcUV5v4ZxOuNHjTsh2eL8b2gm46vq4TX5qmoxGEhl2EUGz
J74QiFqSspGnZP80pbw6+825F87RuUmfKhp6+CJNGVignONv1xagCoYdvNoleydvk+mpyqH2Hc8f
9AOLUhaRiPpogVsBmgxilY4RK9b9Eq1uEx+UEihC9kXjEDDvxwltq/TYFHawjOVFwq53zGT+GqIV
QGoRcB+FHCS/DMJQuN0AN+0DBHoxUtdD4eGL+vktcL1M9txBWKH9CKD1aotJHF/37j3frmRPnjRX
dYeLWKgPXjfOQDOOa+432PkHIWd0fSgsOVhyE2810tVsYl7r9zXNvIAVl9lilQj7WQgJllABm+oP
14YN0/dBnWqMrBcQqlJE71njqWQgggpdV01Oqoz7DBXSE1AzziNrQUjemaIxvZ4bbxYq45Uj2kKh
UjvNtBvSVtMRwqnbxqmRGNTmoBP240Dyw09MZ/zgRwmUXxcblq4N2dYchJ0ZAmkXwICTvnkzBl9l
QylrZz9E5TOWvlLuK/BdINmbGYmUfIvh+pW4xgNte+1ECCHYoJ0IH2CiybVk4nM+KVkcpjndkGcy
eoYF+t+pkJ4dkpx3X1hHPoJSQu8uSiX/Qm1hiz+zMZTF3EBXgJHNlAJEiXiGlhjXNAXseEBojYj+
RvdO5lCW2D+Dg4rJs9z5fUWIigct+cAYziYKT+NxEF002wecPmuim1MBFKMh5feO6zlJs4kA4pm3
nzZUibB3BT0L/dCX0G5IThDE63GJwciMzu4e1/xVXZBZ9bkMa5l+8DcQ9+iextLfY/SCTekRr+QK
JaqcVyLc/35l43CM5cjnPGy0E1fmPFL203IJjLcMa8G/pswOm8kWdttN+6mJEA7sKvFWzRNf23KP
Q75NzBM62SDptFCrH4qRiVGccBRBOp2W+uPnIBIaP5/EXLxbCDYsXD1PC9wfp8rQAK+APtLoauru
48iY3O7PJA3eS0qWM1tU0nAKKq4kXga7SogM5sf6wJD9Fh4IP+5nNYTXi2KCYjAaK2Lj2HNwM75J
N9nVhQyQ7X4Ktc6h4JwTW4a3tQhTIe5NG0xg/fgXlRgPM81F9hJnleMOrijjt1YCEoD2BI4pGVI/
UTuwAQa89v9lUmtDQ+jdaHldBsq1+XCpDawlabpa8KdFHJoWXNFKo6W+YL1rvh+uzKHS1XMCnZln
DBvqNVKlOGD83TEjsb42LSbqF0Xi05atlBKAPUPdsLpqV1WxzrpNWI6c0s2S/qFj/vX7B4uVCZYT
M9JrCZm1glmcN8oKlue91FSQL+KqRPHCU+2zYTxODAMz+Ph0YHWPPIwFprLhezO7+mjHGepp2JHT
WkRqB917iQUyby9DVPctGgInto+JGVuFhxiFJWAPZBmoVKwzr5/mp9WxVCSNcf/qB46Pk9f7weBm
ewTOSbHvPYn8iPzSDf4Jzc5r4QQiWFFNWNDOxvTgel9RN/aAqetKMbdbQbTuUvuYStTg+hO1W3VM
NAbKRaZCGRmCA0ufTXs6rEsB4Z6wwoQQY1cH1/bGWZA4iCVYBzPaQLMPrniIikLX67GBAqbUWRys
mv6H9q6Q7YWKdXthfjNrutsiEfVeuNGnwYtQ92WNLdB1a85kLK/UYBm3iUK5lMyyZqrxK9Kew9GN
GICvHwhCOcql0b0mnJ+uge8PPZZagXEf63WNoeuQHunDzb8YjaIgfAJ4qIt7Ox7/Tk61xVdls9v9
UpkQ4Yyj2Knu4dLFbkFzUncp2pXctxXuJ0FmNgIeI7cSchsVTsXGdjwNVZJE1risMYsEGszJiK+x
5BTgtq6j5tW5+EgTgMF6zukt73fX/lneiObX+3+hLO/jBf3Baq6PjW9O4AIWCUFHky6SmZAqErTn
TkfziKJVjBEUJ1QOkrCFSpnWYi/+WAcULrOra6NC03IBghPzypIMhZgJMTf0JsSPa0zs6A1RWQ/X
A9khuFX9EmVXpYm67I7p6lzY8HNRp4q5I4FzKs3FqstAFO4qc+b/CU42AI48XGI2woLqR2YLUhB5
Pcufcyqi+w7nXfNz1MLrAZuxQwBdRbCR99XX+KNcBoWFeg+TxA5tUYdladb2JBCSzSAPp/OQx1wc
mFp7LrfhiWrl1XYIk1Z9X9r93ot1J7xPMT6r+SJiAwL3p7fku92v8dSvZe0GjIbe+yZN4dwqMx/U
inBLvug1KhyN9mGU+AXXZAGy5++kffoOwictw0dKxHNqp6Ggr2wvsAK0vnmTM9nOXfluuIQuI3Qw
BbHiDzjCwflCBvhe2tqHfr5yIxPGj9UeNdJeI4oAVXqTsP8I9aLbL0D4A2bRT3D6BXjrFBe5rsGM
+SvZy8ERDAgMVNvAWsyAJHHn8FnsH/ZqYm5E5dt9GIoU+SGziov7CEIBVAWUBy6PbLCIkbdWHMLe
NIzLSqBwaImMxogA/KWUhFIqwvnh4c/FyQvz74U6i+FCzUo0WR6MtOsAIdU1HbanzD+mFfZfz/QB
Xkd/14YsTzaoNO3I84d7szceH9GJpnPC4qMYZHMVPHHkSQACfx9JpnNAx4ttiAi2REOq5vNts/a5
X1GJMjf1BRhEU8EqsE3KvWsPQjxt9wH2K+WeGbEfJBVmHOkRj/A43LWpo0RF88SSXBJ26x071nNj
na+a+iVywIYfhvgdGPwLwQ/Px6ED0Z7xZIE8Mj0NWT+XY7dUZ7ebMhOszoSqy2c51dvUVzDLEuoV
Ice9+vbSRxBC0ym48aOHY7nG6beLhKDBIKJfxLiHd7oXjgjwZPO1/MI5ObY4LlV0tmR22a3910FV
EUsktMuen7thiCZdqyzLmgcWsjs96lm28/reyLjAj6WAhSHWr+8gnLRgDDlQp+2X+6jAPmKo2Cjk
tSItRSEj8IsyQLR1jsyGZ4pDvowzeB3SH6kT5JoQT3MOl3usWOrj3TvQjYj07j035B1MrdOdOGxA
mGTC99oqiqnnLUT+JkZ5qTdIOs6xqrgPUMM2Ct2hl3ZNS1uhcqukXpUgm7s+yo2WsPCuLzslT/5A
sVTi2UvkEwnxr0P3TIciVzDfO+Vo3UAjrT6U6yKR8LPaMcn84EjlyYnPT/QAMphUNxCX2WFD7Llf
bzg+R/If9QVBVOyBIYyKMUAX6Zwrb8F6IO+Tz4LOsJEcUEVp96eKXzLPbdilDqYDPcpxh5ZnCoPy
rVoLxr+57RF2lDnulXiUIOj8AxQRlooHhea4ygatzJJXM1QgvC3cvDPtoxV5MhNKQBRfPy3IKgZ0
NFxWza/UKgCOeWwIQHDsOVO0oloSjmBbLd5tAij0LX+r8jnmdTFMx95LgbIji8Y0wqttZpcouy2N
Vs/rkys/u6A/X/eFIZPcht1UmdiJ477Mknn5GLBAXdVDh1ppGr/mPEKdFl8nCz0RXnEbuEXodE6T
xNkdN0QXng3Ksl55c9UOtkYIaauEOHMyNt6JahzHffFk/To2agCEVRk6RubrITZH15mge82IMUdl
Y1za5AqTJbT7+/49wyFsk76pw08GxJV0cbKnjYAcAI1xB5RLBc9wNkQx5MsrXmFiuPKxsZmov1pj
OldoXjy7xHnQWctlyebYUSldzDUhhiAPeA79+DRgwqfWa7WoLtsTqFGLo+3loAO0Q+mCPHCRLz1N
CpjVeycegqOCmpoH7qBHwSbQw3LOTw5aeY8Jw/0f09xbD+tycIP3ynI8e9u1wwCJip8OnJIBIbP4
ua++oBUWrYpt+qkm7UjtaUla+9aRqdKBpNjuFnVRQFhRiZNKbfgPJhgT05zUBpBk2kNdt0yeUfme
HXVls2juar9nsSw/COcoxfYg5Pif7vpUhCpyc5Wq0zjCVRCdrqEP666iuIobuq/DFA/CrQ8x55C9
ABgbWpnvLYiyBHAQAd8Gl0weoiSgfrKzv7uvHvdAzq1kwJwiZIkkykfiv08ZNlbALB6J9JLT4gKb
1xeuURdy7mNJOQf6GSKRR5CPFMs5IgBkvhHcrbMija42/2AYL4KZya0tbZQdkpQBK/kQnzXpJ3jY
4fPIWvNXd79H//fw0Nl2o159Xt/LVbUZcJaceHOGVseN6Qh8KhNxeH0OCdvgBgF87qS3Ip+oZgio
QMeCMq5q35LoU40FIIViX/FNF7eHDPX76pLN8kkgJ1Fdac0zSu2wrPH41q1EK5IfhQ83Sa4sFiPt
+pl/ZslOVAjf6Do4ohWenTEepsi+n2ug3MsmwqhUF9ECe5nnLLhS5IkUph+n9BuE5/FSPV2igFO8
tnis33gYQTC17CYL12iZL03I8RjfoadEaoJ8KYKVCpjgXfW4o0RDEALsioTBHtC7odV3skEfVmwJ
M9l4+XGafDjmUxWHKa/aCZUg+CjYlMEfVd8crZNuQezL9I9RoqdAPdacbbuYQqcBsVfbMvhetBEb
yCv0UWYiTIosvo2ycKh2/5QwWAg0IlAPhNt1VRlCX3pyNrL9a/vhhFBGHwnkq4Ki9dF1MbQRThVv
x+x7cd5SURMpSaudVpXLi4AOdxw4fBtE2SmatrnwZwpgNGSV6NuXsu6kk+5DPtCyp4Z+FsCgUP4P
7N1isJik64JhkN4dvwHi8OyPkwmIPgm0YO4smEaCvPd+Ruyjc9H6xRQDv7BPwPwDsDgR1UaCyvnN
bdr8YLnp6hr1lb2q9sthh7UKe6sjl+/fCXknWV3H4aMhuisIgXxlmQnINoA6g8kUi9iMQOqd5vor
kNG+DPube1Rqg5s/JYXjA6plO70+MlvT07zmSHYJ1eti2ZHXSmCzehPu2i+ztKcldtD1fxlTDMUd
prbcjEiLB7Gn28PaplpN95UWLZwpQUtMbm6LO2/hcSY+f3nJYEEZOzA8IwF2/0DoCA3iyoKk0E4B
ed3HKcq/5sYgDS2e50cFnu8tuGl4IPjDxy7nlHjLAwm3hgDqHH8cz2f7FFQkZvhir9qPFqxsK/A4
/CYT6xHTRC7bf9tRcQVRe2F009+TfYKRQZpxKrtdVm7fgrp/Bow5wiEy211HEuVTKpT3+mnVnl+s
E2a1laK7Ea+sOZ9CWdeJg0HPwjH+9PEu2eyARjCIhdNklc9qB3rhO3NmUcfYdvom6Ou/a4ifratJ
W9b+zA7HGY33nlQ6twISQwMND3M5iTrJ4QgrndAMaA/l6UmUzFOldXA9TZNMJgW3xB9B3KeN0BDn
4rxCpmZJlj5xH+EDctGAZ/0sEkpp7wLNpNJiIhRJWLTXBArQ+fHiAJwLYEP9TF2JMKgEzQvf1mrt
B2vmciTR+92v2clwTJFJH5fQzRZPF2wqZCv9iZWhs17Xt49+OmNlv+U8MSOA1NIQwBgquKZul7GO
olh2ECNPtOI4ySn91Z7JHxbCzXzvoGRU3dF5vbM67rwEx+qEaQMd35W89Gce0Zb5P2kEcmoUlzHC
KFkXQhDxVxbAQexZRQAYrlocKMFWIAoTDjQAYr9ks9vCLHS9tQA6ArzyYzMN4ab6lMUOQGDkjKyG
8B7R7rbA012x5AJB3efaRSbnDZODr3YsfghLtJAdyHAi0ulsEg0HrQzNntH+TEGIN6c1U/RcTKWS
N1J6nQWynYbUR4ich1HbOdnoxncCuPL7o7nEth/6MXVtPHFMtn7FhICmAolzLJzkyaqla/S/1F0B
mgKUQwLBn0Hdlsd2ow==
`protect end_protected
