-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
X9tcu8o4Bq0iE9eptXRhFLIv9Bp2GDj+xa90uLDflRkHbc2CggRnqco8PYzmWZ7PH0AMVwuciFWe
jLQoJWa7qIpGAjchoRzkfx8yzq+wIESiPjgSMFVCyJpdv2Ng9MXnEheXF7MRH7MEutl4TqeWEjK3
q9eq/MBavbx79zbsGI39av4bj8mFtmNqu8fkPe+hqACCGbjt2KT0VNoaOeEZBAWzv2rfFfwQdSFo
fo4W1h8bLx1VAFPOPMxEua2BAt1viq/gtYwEAVPPVnOGcow1egzXSywX5Yn9b8mTqh2Dgd7G+UwS
HKGvWGAhQAoI++GQrWGr6DURhrrtVFQjhoLO0g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
rUCa2YRv9KCKVmY3eOeuXKrc5H7YgHttKCEkyyo41JsgUaPDL6yyJR2oO24yTU2G/wROAXnF7V7S
EEG/2j5bIRjbOdLHmVol761S0C+3As4gfyiSPO0dh4PgEcjK/kwXUkdRyvX7w3qoRBwar/5YiXW7
4fYGSmB8CTpuVdfBpLaLbjqKf3um90gvFwjgbrpQEwFOMxGp4vGgl9Ysz6BYEXOGv0EyOAbOFfbF
PWOriLwiZ7fnJ6TxqJIVk7laKwW8/qJI/AIcs0r85MQDzLpvkTDjwdK1N8T70Oy/jIAlpgH2fCDI
wBBGrDJY7bcKsQj800ajfXmn6YmsDZSA5FdjBzKL5uuR0Upw1zDIzgFO7Rbz9jtB5aSIcKtqnvun
3uD/+zvvMn4p0rAxsFzWhD7dBBfzN1Om2450Nj6sLim16JmidhYopqGKvEdW81ar1r3dLZKxqxYS
teI+KNsIpG3GcIDocXH8gVrk9GOYQd7J19sOKACqBylPW0r0Ye0ztW/s3L8CL5XdvjfEjkgmzK8Z
bxFLxC8YfNvOPGeXirmhY+nfKhyuW8tDHSUvA+mNb+eR+Op8I2w/3jAXYsZrGd4cEY7OtflkbXTy
l1TkOxpU/uvBxVGiEOyDrgIfo4ucYCrQUb2lU85Ars33nDXwebhYIgCO2dGtMV+wCOTXY6TiJ1F2
V6kPUIxtcdN/G0+9Osm4plbf94nOdsZvww2rHAAKmrJSwPfwpg8sJRH/HjcIo4Lw+Ya3UfkoFOAn
JlG8AZbXqtFsX59qPWAWGVrvcfMT4DTU9Ukohtr9FLZSrqhVmN9FWCoFqK6OeE5pVXHfhknu4TRY
2GC2QyDpXMluB6I87+bUnZQGfYJolZSIAYYFTI6EOouFwFI1CV1zV2QGxq20ay1oPn5a0NUjzdX7
VKL5Ycov5x4REj/YqVOvNO2HidlX/3sKiRhmB45nW+R4M0T5+AkaJNYaOm1mGeXK2QMf4dKDAT4A
zkgKZYHvEwAvODFjCIkAA6nxuTX9cxsqK1/HNpTL67zLQDkdG8tnIwzgBn1xahynzKdx9uHljGxZ
4rNZOx29nAbcFaiwCg2lazg6UoRFDz3Jk3XJA86ce3vMFmSSbdj8pF7Wopally+JGhxCj0Tt1fUh
qCBkanLkHZqyByzmj+s7c/slFuUFwk1VQ1MsaNuRCMGQG312LMst2D21yg3XxJQG7fjKPdkxHxB3
Joa3C663j0mXkVivEqmoAgfqJNeuiH4wVAWB3fVRtIQ1xk4TnqccJCja7p5qCXB8y563YPINI1UL
fz2V8kP5V/6C/EPnEqDCL10B62KvM9sgFZLxDOnTrFe7G7sAPgMAB0nu4IGgptmsEYjAt310ji97
ClI5pRba/XW8KCYjeKso9OpLaULwUiP3XqBc71Edo22McnhfkjY5HLFgIY5v4m+PxGKA2dCU+CkO
Futvw0QEmeidy/35WQI/r12A8FHx39iMTJBrvSE3tNU7E4/QEDm3EuBk3JuerJmJ87WPe5i1kRzK
7pWfjluhO5T0raFj6sdf6vTzVvNS8SqcNOIoJ0PBdRkMMPGmXfK7bXTK3qoExY3ytyDZhu6kD0jx
+peaKXxeXivqBl4+W2gCYguEuGcDQrRgu2I0wV7NikFQcHWBhZPPLSDIoAPIsVRKoKRKgH0A4Sfj
yYOmsuAnR9RJOyAgMvWKLU9MIEgHwm7vgTLv1YLBQe+sXG2tmX93WPZW27oGbStK/nGUKDFxwKwV
ndR7BGBwfbxScvtmzU5NUii3JkidOh6C1+Xl+yDgqBRNYz0W5tVLsMd68koi5WdF3oRQmzk8M7HV
vBf2xU9xani4UHOhO7tq477TUsAig/YBiGJcd4nLsNpeYcIOM04lqCfqZj8R2mwQUUUUqvhNYlZJ
jTItuZx7z+7a+ILs5S6Wk6MtKQ4ofiV4vgpalCPZM5DoBY43d7GkINb4shI+XHwaWZGmxvmqkSIG
V/vlyFWgnudbmI3AGCqXnSYsXqdrkji83Jj/W97xGXP/m4EikyZzswP0qf1kNGuoK7iVETclGkQM
iKrcs25NMqJj0xWcBahqzF7nqr2hXCOYscISkR2QoFzEd9IoTjJEx9RXGnxee7t0aeK730rGy/kO
4LgBtNSTF3FV979UH762+q5orrBFaBDTeOtS1MSYIZ5R/41kBvuHQQEMqTK9APpJ+5bC/Q7Unb2J
MAoYFJkCu5bc5ko59aS1Jnx7KoYGOn6o2LdjCHZOR4COlhoNLTUII1Xwe/Q/Hsxjk9lZbDcc6b64
hZYKT20miJgY5DuisJgPmFZikvifVI/bAHRINrTaE4lQEPRryai/WjwhCHx95ourg33sKYGmOlLU
OmRC+2bukOcqz/WeFyvUj4jQD/mRAyurTx7Xm5JSHo8gokAzDc5BgHvol7mgKC86Dk4/ebLxVJ1P
1aHYR7lohb9xJKfieI/BJ+lBva8munv46atrWk+tF168DtBGcw79Ha+3E8/A5alpXcE2gN0FWTlM
s7K7Egc63xrE/Q4QK+w7csugxnU6w+syKUJWD1tEnfdYCPn00Q75H5ZnvO5kVLGaHrs0alq/bJKF
8YCnsqRV6xhlrmi476jOj1IlwT9xTRUkJu8x57Kai8VKsUP8Q/6RPfZGuqrm1EcTiw2F36BbG1II
ZgLdKT3KhwvUWOcntUnEIkpdTAqsK3NaWKViwX/IoZl/z/d0XjsR6yyoLYI3F6ARsG5DlB9BSD+P
fX5wSlGRzcRjbOOWqa2Oc+RSsrnRtBTr/Y0m7UqpPFnBViducYveHZD35D2iV4yY3dScJLItBds2
t3kz9rKoLkUxgtAylbDYmTjDKmdp0rzTxrw3Bd1l5IHV9iQhnQXs4acRw6Um/z5IcKZxPSlPFH1J
l6hYSkRckgm8+u3NTOkbf4kTX1MZc33q8XjchcRVftqW2eVvBsQacMAoy4FY/hpUH4ssTfiFOk4I
o6NiHb7WAlvNXNlspO+278UW9FpuvhNlg3fQNEXXI4bIBLbPrYcyZ7kxAGW4IKyHZOqQL+psSuWM
tybeJjgqsM0+s6r0n2dysfMmykHmxnERCzjftWr0wrO0zCzGRHhYYUkHhMGPZJwmhK/J3B88620K
owpk27Ao1bU/8WYUyaUoXm3VuRSuUvO2lLvbzUhW/zy8qd6lvCL57R7cZHSBdBgtQPQ9Xmnvqdkn
IsPIpuqdC1DPsgAXIj2DsxD4/f2ZBT2uGhPuTO8K4yNfDtmFC0JsmPvCUeZeHw/2T/4BR4yeJJ37
Dz9z1ZzEH/MBRViJpn7xElG8irzw+DaK8Jq9PIjMPm4nzBXi8Px0yDH8ZI6uCj61pXsJ4qxLaPgo
57RwuwmPzdItQO46dvRBDQekcVqF1OMBlVZ/aSOfrxHgGl5wPx5IkeSFxVu6CdnX6ALpzLskhlo9
PQvCRtBRm6PqBppZW25RirrL3UPpXrH7wcvTRN9PM6P7CoqvB9IQrFhSfiHQ81Z4GyI3XYXAM4YM
EYfzj6bMpRueK2Guxc+WOq4tXrM2KjXiIXzBudvE8gfIqDa/1Vb1WRVExbKBoS6psD3RGFKRa+8m
YdvSN6JMYabh6rw7n5vtcdUA8iW4QBI8D2VjkCKQ8/XvsZAYBSofs4ibXeDUhc7KRaOnX15jL6Tc
BPyJTIy3fsHVHqGILxNKZ6ZoS4Umr6Wj4UlEmgAgyZ+RqOHJ3+q0Kq/UEOU0j1IcfdaLAuOMqZVa
aPlfC/zG0K7XogwsP6G9xh1CJEfdlIUu4wQEXinA0zWewGLEqMgA/ZoLl8lOsNxN95QVQycwNs8I
fP9JQ3k9/i7sBQ6nUX7AdbMf8SxazpLd8NeAdLzf5IEy9RXpRU/JVM5MnpQZ4pJZQsaBGL1+dTdQ
lP7bAzp+uD8C4gTk5bnk16jpRE8mQ+q0w7NWjcE8DwCMjnEsyFgUjcQ3dCTGxZiXXVHKh37gzPnO
RD0rPHJjkr/e+6L5ICr3S45rY2QyXw6vNegUPE0cY/aVzwqI8B9s7qamrDmscdMpYBdCPYtlp+SO
NPhm1jR7kGkaPsUywhdthwjLB9jyiamKZeMmuVE9ppyJrYJka3i2lTZUfbjBsVVOoJRGt574ZeHw
39GKI9cQwhUXMnG0zyLdxpwZjEC41rb/KGX4SVcEtpPXz2ScI62wz98dhQTxzJkTqpLuOSGSix5o
7E6bOK2ZId9eeiUfBPldNaNhcnRRhppNeJrGqwcCmwhtpaLHlb00lKT1g7w9Z2yTApe5HIH1t5Ju
VreULO5wJHJe50GL12yWdK2HDlAE7Og5ZAExP0lL8ZTtKDB2ho3gqnfNnMdyhEiKc5SEYQ4v2033
Hx6L3Z8PSYMHckKQ0dl5WtTSUWaDClVgsHBWV32L0R9+bXN64wYeuBtOLL3qExJwRzsKDttSF7MV
VVafP6Nja+ludYvmUsmHaLapTEZEFT2QF28TNJdGEPjnlF5bJ8JtCKjqpTmq6Gx05DWiGTNAk9cq
uMO5r1b7z0ePWKUi9yamfEUuOBZh7JEjcGHjqmAFDSuD8V50rFxhBpa4wl9olOTO2HfW9SLH7nPh
cSrdqUDBcjB5Ln1VOUjOZTeYvbRxFPgIW1ttL+kd69hZgFvpHlMB/y9CHDJtKkLzOrqNPiaHf2UV
ZmIEHflRI4RXZhYBV49XW1i+sCoDxEQjLPjrF5Y2EgD/WjZVB5ihdq3UiglDOtpHYSAmfg7waSPH
vrGDx1yIwt8BJ+9Ur1/5uYb2oszUbJ/zuwC13rW1Zy9l90OT0LVSqRvI+mb7dVBIoxv0sPZS7odR
8R+/rS0EDEqt2muRfZMx4cxm9kEtVRyJvMDZ3ThkD6oIS8W+eoqAWuGyPI7Um8q0py1pZ4tb40qk
XT/hix24xqymgBBrJHhRee0bIq7Kf9lEm1NmpN7I2HYr0DQ6nkDl+4z+CtN4ABPh2oC/aO0xnyZL
os37iMEoCgLzU5Aag490ROHMHLxKZOLDQdcyVfCLS+Cy0JX2rKc/5qwnxyyW07Ns25hUYY/JBk2e
L1YYAEDGS/7SHQEaTP2RL0u4FjaTJOA5Uvz0y2eDg1Z73aMZ6pLE6VplTqho4REgelKAg7zyLC5L
xeMyGvFMm4PxGL0Ggl96JCg8S3E7KNCYgXelOItPHgSp94nBLq/GgxT8m7SiB9CUXFJPcrds4Z1j
hCCiIkwX/cK3fIPYQGZP6uPulU5gdPV1acBD5Dw7RyqF0aA5Fm7jw6UrR21g2+GADf1RpuoxO6ck
c107kLjRcD4LfJtG+4pMJR0cwBH1ksMILffZ8lK1165VOGKxQZfNxYA4FrzFcos465yadCXWbrbR
uUUBKqx1EM2D+HA+Rptanv02mL+LIq8QJpHmTjzO91GNmZHk/qyU6kal9RuHXGFALROThKFAJZIC
8dHD7ojQyPVoMRwip7eJC0z2RX2JO0zLudYS1/Fa6V13Emi0m6dhSJYUuteWTaYZn93o/nj8qezp
VoQEZPMXiIfojp4bwoVIql+7cmU/yH2uSCilTpH38fus3GgXjNA5y4AbH6nUKIt2gM+0SFasydmf
XTcU7HGitG5+KzChChDvQDfdQ9TorOjnEPKjDcSjfUo0rxAyIdXT4l32QhU3IWomqGmTOj9vMdBd
ykSObDzrRJW9MMa4gqKI8og5upOLi+IrESK2LSHHL6pClmsA+OdfPgPEDvJiBb1TS5hH2vUZd5OV
Vo1KA0BYkjT63lY/MBaybIGgpjSh3wWdtZvMaqv2KKz9PcpVeWj0UdY0TQqFml/vXfKBaqCiBtVe
egDYFvbiMFvfLJn0WuXQ5okKpZOWnUnwpunhE0UIr2ByU6e7hFPZuaggIGyoYrBet3lKycz0Yte+
CQ778YmRLtQWYBX+o0ffbfHzKJkaKel1rhvgfWi0MPC2y0rMejwHazhSBLih6VLsq06LJzrGfo6F
H7R9KXwplVPg+F7Rp9H/DqjapkL3DhH5SdkeSPTRnz6PpYn6ukYGD9Z5qz4+sGClFTamGaXcALmo
17QTMjJTNEMGnNyYFTOBljj4stq1qMLWo7ViETxIK2YMTt+gqA2P/gHSm6oj5oWm6l03GYpqpIih
zYXg7wTBzafku85D/sMG29Gv4Rg8QAWaCJzg0L1LGGxjq2OjNAqbO/TwEtb+8023fB+0tBCVcylR
HOTq2egqsQaLN4ijiDWGfZaD+CBa/f8duhhCQKjRjKQ9ZgGuW4v0u9fVO0ll/X9F16MQgYgCYWmA
a5OzXEbJ30rg2vHZdXr3K3KMq4OK3xC0rF30f9etnQA2TQKHSjG3XaMzX5AcXPGLfCpwsxwVu8oo
PlpnQ8IO6nJunZgkZb2LNVap3xqZxeJ/vcGzdwmc2qGrDHGKSK+hFgv07Qyhzyfa94GJi5gMyFym
0NgkfIZ2mtn5o30D2e3161b4H9SAtSLVpmtVeZZzXABACqPxRhiWpRIcNsJU6vuLTI3QSMdCZFjI
+1eMBmxyvXC71hVcQ0qhucoeJ0xP2m1ZvR6Mtfu3UO5gfTLXIDamR/IB/1K7OO+F5qDiu+V89Hfv
VhrEXOtmA5spKYyxIOrTojjkaO0eKxqUQSQfi44lyPIR9iJnddELVhn4RQC85IvRj6YKrb8V9ciy
Nbd9MgdroaParGOywjt1mxc1fiSwGUBONdwV4gfzSDYaza6lVoszXPL1aWv23b7lKh2DMmAr1OgF
WBmOkeC//omw4pQH2V2EDMac1SthpjDPoxZXFd+siWyQpDdOxz4FdO/zAuLd1YoY+sYjBIATQ+6/
vg/qEWUpig11oOhqncOHH0A1SJBdC+lwOcJ6m9snHPruCNuup19wY6wUiUtMHGtpqRCzRIGltVa/
59hIY4A9kUP22+8yNSC5TUATKgw/YWK45x0NBJZd9o0nCIA++lWvVE0MLcanaqosDFeRvnpuhePx
95w6pCc4zTveC5M742uDzXEMr+aARYHbJ6h+Z0mTDu8NgBIkW5tzRWhOt3F7bK/iwDKAagE0KoG+
kvZfYCRp9Uti2PaQQpoS9VhM/43VnzA/f5VIcTHUiSBs+D2LM+sHDwXrA05YN5f0SPTF4Xejtj5w
WR8cp8iiUgf5Nhx60dJxBGWSpN6eDc1XsZAau91uvKJHjNbj2NGxmWeDvpaJfFgdzCgJR5qmgQV5
uuiWkx2ALRVAafHn/4g9H5TsFBz3KlC0tp2DV8ayG0VDNkLEZZcLbX4rihM6RHUAUoeAcdIzxSe8
FDd5xH8TnuKLEuvDowgk0uMqqj9F9f1aR+n6MqicdMK3SFv3sy2QUkJkPE7LSrsF7e/MbK+aiKIV
o7iIZjUKmXEZWt6VncznQS0K0sHxFmXdr0gGaRJFXQwqELkkWMxH1UrCI1ks5pjsGYKAHH0FzYFS
Ljxc3cS5aFEjPrOLEbafji8Mlpktf2thTVnNvJQfqGj75xWbVgMDw8D22AGOauc6VfTqkOMsZ2c9
FXT0R++770RDuG3K4pbpzYrP67fkUsjKy1LdNowL1c72PUTFzLZ4P+MmubW32KxQD/U8RW0IpHq3
R9+2bPZ82gV+Dz9KD9TkH6JqVVN7DpnSsuKw8J+GcXRCulBXRvLR+BU5Q1aEmKnEgj1Ru5H/FXlo
X2KfA2sdhDnkyZdN3NYGkoogOr0Kg3IwLeFVyMknkaHgRQ3W6HCtf/UrWSyQz4aJYD21ZjyzhtNs
lCdDj6yR9GnmOTrtALje8rWGYaQkktWm3R5GFhxwp3XJ0Ro9BBADAinBROhTfA8ygIPNzWTtRFo2
cb41GX6AaDJO+O9hG5aOvTXWEa+Hle6H776bWYScUYr1MkE/3VYD1aj91ZOdj3B6+n+rgHMclBja
mHHYhI3P6pJ0QzCUyfNkL3Yg17M5aljdNbTDpnsFmqmz/nSklJDIjD6DhHnjJjcUeF66yPivzcJd
Y9pt0g6b6RhosQ+E0+HcZrdYFF5ayhsDI5V7C1r50nfU73Z8Age8NC2MQYsZJVRmjtsoO2J3sMeq
MLrAWqUhxV4KGXoAfZN7hFQZUGgQSWBPZCuHbz7cJH/Tz4cAJWBSS9SXv+WGcCqQIoY2evpIanCl
lFzzzB1xYNx/bX77tTrIgBp3EL2AOkKxDcSzYSCneXrd/qKmARJRa3uLBHTf3JLSzpPPwrrRPY5j
z+X3LycCEvXMg2I1ACb9C4os1g5KWqlnjFMhplr5Yeu980eKj+1doVcK07hdybBWpTNM1B+jL+r1
UaE6/UqwjYiiwweIaI1HHZzep/okp14g9kvY4GGeysp6Bc5ctOXCqXNhIuA87H7DUTR4R8PvIyMV
z4XY2KvZJmMQg8akRfOiOAVHgOslcerwZqle2djcJAYYkwGc3nXk58yfXEvGrq1bvfNBRUNiwo4U
NRtF3LTevPZWQFFu9bo8sIshGYmrM6Zl244DCLD2eP/WN174KjGeIWKSs5MM6jnS9YgtbNWOnC3A
8/AZpxW/o42+ACLJxVhW3MROjnWr/s7G7E+30XPAF4U3frcIw56xbHoBhaSiD0RDHgPTdWeNfMnx
3qVi9IEjPKtE4FS24aN02UFs5GnAtn1SqbjtSD6uSXqH3KeB35StpdGJ4B6e9Mts/yXp6LvFTc7Z
Dq/f/2PbZVFok7IMz8PpgIv1SJYVzvcF+k+ZIMM8kEynOmE4qF0/98FDQFRYFLWsoPdi3sZOA6/Y
sry+uTddTUXtBqBMvE9lWxfv2WAPrBTyU9TM8bN/HgU2DzA+efDwt025VVEBaPQ8otqGJRxHixaU
e96GwGDkS4caFYY6c7iTl5jSnZgInCm7/UNlY/wzLro8g26/WdzX+7u/jktMMgPyrXStvXoqdKWz
26G96m6VTFpo8BaKPD6HH6PuIb44f306imFtoYfGkqnM/VHsQtIyyp/tPacD4vNE9R5jvkMxrykj
tbaT0+ZCuqMbqNuaM/HxOpUq8ISGTj/KwfwbrqCq4tZjCzbwfYrxV4pjTOCFb0pwLe+mOFQpnH2y
uGwXQUl+LNUz2NKGrDay5olTbF+At0gn6VBx0aDZkTFfLTDoxhIv1mLz4vgUrVY84WN1KJoPElGP
zujk9pEzgr7QqNgk4Li8g63VE0zGMCsRJJiKxkBjteKvMqIjcuqYMWv2UCbS4vHyqc4VQc8Wjjyl
EaAkq315UHYgxxzYSiDy8uMMH5/r0Tu4/8/16ELXYGl7ZwK/J7eoyiGpAIxE0PdfBl+wUdxQuFPZ
Pvbu4y8u6xVIaJWAzbfhCEb6S5CmkwWLEf145Bd39QL++PY6zwOtL+cY68GUnth0kgEwfKwNxycj
mfcyznwZpSmqrDCKza0hcxQ4iDRUbL7tXCbAdJ+SlIvPIPrhhi5R9onbkndH0yJmd+gq9Mt/4lhZ
7vuECTsBOrPeUbRj5ZooIdEVpR12fCOgvY5wiH/lBFg46YxbfrUMBSWgPcf6Dn8XOJj0/f5NCqmC
qmnTPW1SbQWD4gbzv2lV7O1w5gWJccZK8/+W1sfE9XQYX3aU30jmTxsITaEe6f6PxYeZu/RqChyB
MpxBp7TLsgkTt5gcy5gwsxOUn8KjT54RdjpBffvM3w1pYSmYyz/+z/OQCUnb2yDP/TIYZJ6TxIlg
XMH91bzyaXnViQGUSQtXspv6iJNLrPopZ7umMPRIPyEeZPXTC2bUgaky2UwJXOBd+tjoWOjYskH4
CZYG0lppZkJ0X55EEOOb3U0W08cfE46yZimUPvw0s06QBG1M439YZs2GK1ggM9QbACUe7cahguXD
znMMMyQYhT3vZkLeSNIgWhCRV1aNIQ/0VHdVxgUKGio9SshTsU/EJdUWAWNzcUwt+N9QGT2W5FLJ
WSqV24yBYsxPIhAwy+xfMfZ+QnnMxjDbll014ENEBQxpjtuMM6J4pl8RHRGZKP71MJgXlAziZ1Lx
XsLbXMAAG+RM83GsKaEww+4ymKlGIgPQVf3dHN5cfQlWuauukqyZFc/WqMGjsCMvMR9MgRCE4U5c
/44XKuhzCGVC7oo45/kVFrd8rIkskAOYjTdc/b2gei+f8fAT0a0LOuXu05OMo9PuvKrzpBbbOinB
mrHyXNkQ3uioxyfb08OSYHfdOW36c+kBgwICRg0QN5BnY3UMAuM6Sz0dBpcHjkvhBxEnDEhPz7Xb
m/yK669erES3D2r93Z6fOb7WYoUK0MrAnHli9gbXCgxGN2PthkqZy4J7HopiSwgg+ufK6z+83WF1
n2J7Np2DMTXhxxBOpoi3hGtSs//D4sGqASH9o6T7TgY5WAqKRozWW+F8nxiKxBXCI/oLeaCAisXS
JRUbtfz6pEnwLCq9wNIYywKOLawbzHVKAFk71NNpLC75wHr2YLa/GJcdEqiVt0HgcgPmrnZDhqXl
kVUk+v7o3bH6aMsu3jdg4PmSQ9/RGGU6hVxWXbpc/Xapmt4lR0cAKA+lgJvmsrgZjdPhg2oXqZ7F
I5AkRAlRDkBu+n2KcQ9ZegFwlCnPrGLJDawfOC25JQo3Fcefq6qDMRV8KpxHOuMUYl2wdrATlidx
Ug0p00Ff6+kxGdv7MsS6qmJtN9WimvCOhP53C/rNI+83NzHKTUww50fBtmljGArWXRsvIa4xv/IH
5RuEnv9jWcxML8ZCW+VyXqDdYbZyXHNcoIwBOQ8cnzEzzAdZHvHbhgaqlm5+boWl3V7jvOlJrIfW
6NDkzHZKrgost092yvr0XbkBRMOWpH+whsKYBxersmeC4t0LY3v/j69JxKnPPgv9PnYH/9e1NWdV
BjAcf3kwGljcnL8RA6m523C2j4RRUytWVdCVJn+o/0A3hWGTviPwy0flPZftYN4VWrQWFy1seC/W
EOgbA1mBO1Sd4aZ8SeMUThO5cz8sZwz/1RRehDptOJs0AWHFBbe3O3kgcT8BF3Xi2C4nwTMQRwna
Pqhl8GFH7Noi4FgxlyCiTFPOfdG0sgJK/Nv566y6cpf5VAs7ZPzhPVj7mGMcHs8lykbI+9sTi+mn
xgFUsZEgCKCydaNI6AmKgkksvnN45B6FyhdopO4h8S3VvBox8i16d/KOTBzg42u7KcwORYI/dgyy
Wf5ArUg/Mxjgk43Z3LroR41j0NpEmYXvFECHzaKRvbDKeuHk+92EVuGRf6NNkaXfOnWCGOzz+Ukz
rIc5yVf0bNn5EQgMrHl6oqi/glKmR8sQQUNuedhXD1sPem1EXYiHY8WWkb1DkGPAD9m84x2WFyYo
hHJZrBU+USE9wiv7jkHvJSed70dt/92j/gfGDRIzxxhwrk4U+012MiQCrLENZfAFWMjJ2NB+K2fY
YJVYDMnQ72WvYiUF4IHQyFcNaId0SHqrNSCf+7gY32tN7KCXThQ6i8F1kgewEO40spYqkpWmE2q9
xbFh5TB3/Z8gSdDuiwPfgKqZPQH2pNhE3wUkpk9tACw+kVyaPML+SZvvWIAZCym1YqUwtTgwzRXT
ItnOExHW5nqFiJYM674tM4LsQfjnCyiMqmHGMFuNDiqhVjlIY8Yq3j43/xu4crJ/TaH+H4RjXSLh
dgNgzukfbtct9MVF3hEEAqnd4unYIKbueoceJnDB0YAux12FLwayyf0AucA1cbTEkh8Nqxb97s4J
PbVRU0omkxc5RzkIHe0LC2zDg66Bjp6AMbTjkSRCw6BqAm5cO/pD0opRl0oNd6RSVRjcRF0phCUT
B834BBSVNjjxZcdC5S97n48mtR4Lmme7KFvcxoBGbYBUsduQ/JmK38VvNYjuSuCq+gXGO7UiqD6i
oJdruiGb1f2FYyytXMLMFBBthriVrAVuhlhZ9qdQC599QNyjbrb9SL88Va0M0DKBO2Nr7cI3ptB1
miy0/qlB9p8kCseTN46kUJgGP+lywEhR+39yPGAfxjo4T8qvjNHVptfjCqij/sJNOyjzC6hsOieB
J5aAeIGxG5Yd8mrunYIn/GWCINIG+DZPc+Oz0oM37X6S0AuAS6uIBiWPDceX8Dr5AI/ASsHGvDJe
KybZsrqbO7fXsFLTiTYux76QPj9wacaTFggd8lD8igKuOBzSlNS4gEqC0bisTsH/E7AxljiqPvaP
3XNJWPtfy8kAsuCUb8rvjw9Du41L1+w4+JW6GRf+CV419ws2+DFEkEVxm/KZF/fP7hYrLf1rwymG
KLt4mdyIgsgJeI6DOseOXAXzAt2OaId7X2R3lZrBGGBDkHIwissgoalXND3N4po9cTEHNeFxsoSy
EyQwcuMbV3cZbb4f9qOlWNmIm9W+DFIeM5MjmRqz5JH7REBJBKKUHgQ6Jd0yFLjW7jnoIJArE0k2
dAYWQlHZczHuWp8hfmGHXKG8NyhBZZ/lX6hyD8Q3EtHt1ClFD/oZ5erW8KxKqma6N1TScxY69JJF
3n6jBrJFzJwEBKoQUz3jWLodVXMMOELG6zUZX9n/hIDBVcK2OfrVtBGLu+reKzBt8mBjc4s+QnkZ
nTp3pqiWWlZloByaKiGG4BF6wxPXG91hpvqQi8QUPI6NAiAPV+Gp7EMtNQWjmI9aWnT5RCYuY6ZG
8IZooIa7/EMEUI4BPiO51m33xOqdjezq6nApSQM1a0s8lw/Rn5qVcthEYKCpwPJbHXWasHcgErwT
nM+FDShFc5rXUEdTCWhgSSTHoHNMDskuTRPbmzdm6XjJpt7zHdduChy8kM9w5Mt6Gex3Bg/jZnq8
5J+rtVHJMxzjvLAp/ODv04OjYBAV0cB30ahKU3QCWc6hUUFT+Ua2SmOUzFw2SZO+gA/YPs6wGjKQ
hUyny8juvyKJL4cWRZTGlDvLiNphg1c1nnz5sArWJKo4Di8gFPcct6ZeA1pmyyQ5V/I/UIh3sJ75
bCDX0s//3HD1Dlmnhj7MYwwuG5ZDOkTLiyNiEmz7SEHI0VB2UZi7nV0F3F9SkF3j2zCG7SK/cSyK
R36AayDD1p79BEejId2Zybs+D1WC8Hq8XQqoRi8tJKZqwZwy1nxjGmsg6FpufeCGrWFh3lor3dk/
zNNGP2auklnM3qB/RxGcweQ5FY0zt1/yC3RC0qly1WSdE3hgaX5yxgpK4EXS++Ed2ytWavTUQ12R
jLtnYunuBX30A6mF9bKJUfMLUF4WRuUIPosWr4ErnuZpFUtVL6zz+1khZfDy1A2VFZZ9UubDkwhG
moJ0+AfyCPPiBxtxBwS8HLobv//4lXeVBgJ524BI0KbEejhZgWyKHr0hjJOJC2uQZzKCxNufLXgP
2MLMgI0IwceTDP0UvVmBtCQdDUQVZBkYY0Gn4X6aHDD6ZqGAmid/+EXJGYJ/UHS3qN3mFrCmYD/k
73VUaIBsFvUzJNuaiCx34f6ZRpyuF6L7eYPsYtVDbAjUNMwMWae3+gbw9ez0SJS1F5b29+Fqw0Dd
p70Hacmpy5XNuscoBwnzz9zZn71g2LhsjJJiI3KQj74v5U8HIXO1jlCHcMwlQsepLKyWzr/ZnjZu
CnTIMmeEEpwlbwI+H/uLYZT+B1V9eS3I28HVY2FYUfAJVQWsx/5mq1lsnqkcY73z+B242oRzvy22
CPYuNZJnZMvp85V7mcUikMJ75zEDKJqM+tacQ9XNd679sKPb2N12sgSnJ4LrBfhY3DvFl1YHNnIn
+IdWCy+AYAic/WsEaJ1gwKcS1rrQLYHEvnhp/oRlEf9lK2WVUtemoMzW6w9E1SSsuZsObUh7BFlO
/keTTM74HxesmZ1yEnBdeNHtWWr7sZmGaIsa4kuhAdOj1pBV+m+vI8L00pDw/QE/VN6oCa9e7IRv
JDDWNouKEGD3Jw/xhDZCRWpTLZbY2WsEtilRXLHKAQTzDZx9J0Y+ywTUVuRE9Jb98xSwhY7uFmsq
tiiPCbrE9WazEv1Vb3m5PT2mVksGhNzYvTgJTfprVoDkCTf5jtdkqrW+IJfRfWniZEzR0k8+sR41
7zOXPa9FMNq8Vc+jqxXt0myYSx+JnNkFabhahGCfgEq3JZXJwFzT3hjbOoTq8QupwTlkMzcXM+Ty
o6TXoPviqJVOOjO4LLFo+UPoAsExILx1IWdB06ored1P7BT34vq/YmhErCukCuO3vuoJPaPk1k7M
s72lDDDSPeZYkQN6VRRLjZGr996/WKV62d/dJ0bMGsMD+wbU+al3R6JOyYYjDsoBPgjuV9eRG+Gj
jIF0yzF9bHv7EqMZRB53kogPbtgkomFO9DLF41WrQKA97IUGpK8D/iuQKzdK6OYOzXiJxlfusy38
HAvtyzCrnLL/ms7b/3n25IeIIXxLuQXs3uMY7OxIPFP/59s2YWwDrSTDvwcghgJtfK8iyDUr2aFn
P6JYoqhe5WRj4eScQNOnnzfddhbrLWkVi/3lc103q5I2LANb+jjBe2AQa+cB0wVjA6jpQV5mUtfO
l22cNSyF8LetOlI9g3OP47QIglFGFPK+zw6S8uUyFmsF5E0lmoM6+tDM+HMOZ1K5QCYS+MIP6LTI
UIMDx+g4zp/EDhT/iYRxC4CQGGwQTIh5y7Vdk5QPBdFnqft05ijJ5bqBxa/EHAlYhrWMbv+H0kY4
zfs864rkZoiR96HNlB/AQi9H0oYu0puco+AufH7Tnsj4obYQauHT6a7JnOeWzbRNiBnwLnXJvh3t
7qL1RiMiiiOzFmbZojnlJW+DwIYpkA/6TqS8kmFmsfSBPb9RRnUFnTcAS+CVBlu1ysoN1DpE/C7s
ebrYZcy8Unze/kuB/Rr8IrSinKf8OXihZUQfpz2xNBsnmo6L+uKG1GSlpo7SRjj8m/sJYOqwEBrT
OQQmYkDeEYIqaZHFIRQ/HUAKjgPUVTYj6v0ptNu0lEVthbNwVblYmXiCeLw5qaDAcC5rbHIWZJPa
X+2nRwneOnjzQeoBEHqNAeMozWPYDw1eF16wZ5fQV8btUcGs/152hGxpqvETt0Ps/kjr+K9sMtSR
uqNmngwJGj2e6ZsFXDRtXdr8wWO18kdrYKrXcAHrZXqzp66I4hJDGQTAQvCBO2gdwA6YM1VufBrx
J6uoFNJ8vsfvjZ1OAxhRpimIHUEeUxccikdIEOFBP9IaqqglNHZVxg4SqCICwtssE/6s5/rbFi4R
F3pt+uCbl5q0APe8xIm/Erb9ybhbR4m2An9wVYUH4sK47ewEu7XTfuBKRI7hfuT8Pu/JTkRUCFKE
cpgVOrsBGN6PUKjDmpX9Ess2nUMn1FnhmlY8U8DfLw+U43vA7Di6HE9GBlnuWZPaZ93HCXLg4pBW
omQSJZ1cZB8M71+evPe4zdBr9VW/qMtlxpZxfT9cmHelRGicI7lGTpukogS1Syq+Rtjzo8EdqtOZ
DM8xX9RM/UWNV7n+AzvdFEtdNwZ7Nhqssxygp0E6cQ+IwBsbg5G1J+G7mtjjDnqJC7y12+BbqlIv
sKP3iOJ25Y/TIrIqEUOEk/auGn1OEruVYHLTfryxJLLnFqAdYgh3AbCs+8RD+8l0dTVuOG64qjfw
ecD17QJCji1ddSGkmasiEzF6b8oAvaqbcwy+8GmGcy46oEqtzuY6n3sRq+w07+74pcYvusapxt71
WQnjvFZU38Qi25h5kFj1xronAz2T4oM0RFbZwEWpLX9xRUnzM28/3pJErVmBmgbme8P1njgOK8uO
SlpzTwNw7KqSE7SvZj6s5IArbM4lAijuXLY3HX8Dns+AbtKcDtz7cKqFlBrKeYYpD/wE29tyayvD
S8iyl0+7+og0JaoYYpI4VzS4oGPopv/zQkxlNjrfmYZvp26efste3T+4m2FXsZIMm9RpySRGYTyL
len33xhlEVuaBXzegqZZK75TZarmOCyp5CAzrX4SmmUVlYvBXU5Y1460hT+HERLfaTWnf3xWJqcu
/PW0pq7hPrlGVb8jR1iNVC/kHwXcibZNrDP4iE7FAhkXJvJNDuevxqN4qOfb04KCGsrVmsAvNMS5
eHNJVXpA37qprBjfMI71WttkujYEtLMqCZJ+7TvkO4LREDiuqgv7wIeUdkMMNbA16tMaH3krhweA
9RpnqMEE6j+ow3pJeHE9LPXnaXISSH2pxzKli5sY+VDpxQUrA47m53oK30W0C2gY2FdQcGZlPl9m
GfK8KaLWQblMWw29RBxtEjdheZX0Q80MP//VX+LVtVDAM9VzphLm+VEjwfMJesvwigMrOv0H03nD
mpSY3aZxA/AT87qNofDXrRzErs6aplymrpbtMkZ0otf1sJSAOxunKi/sQvgpX9a2S75lDO/JkRWk
pZKfSpMZTbmnjwu3laiUeV+da3UNkc1lzVbBCY3u0mGTjmCZ8BM6KyJVTa8HIqu0wdDmAL565hwX
0nCKbsaUXfwn9GE8CobE0jSptf9bx/ptDD5U3ioa7WZ6UAEr8YKF75UuJXhIavBA96K2tn3MZXWn
DJnfHNjo2CIz2dJzeSpJqFyOell0FyZoiRIhoORBQCnt//fNlAWyfJLx0FroCD0xnqS40Ivch6R/
nRC6E1EV7H//BpiM1obFQvE+3/bT8piyFNN1fAZVJYium+GGWBJ+m0imPqO/mWEEMGW7OPnpkObc
sH/0l5o+J7Q5sUNnDLCqXF7IhW5TEUnoCV1I91DZ/SVYQLrQg4Sdl/4bWwCCV5QSvd2WGA5oceby
HuodTcfoO4DVRfuX/U3CBPglPZSM/kaoJqoAfWZcP93hXOvUekPR/NajxkfoWfqVHg4sy6g64fXJ
/vYQvE0oJlERWmk3bzBzLKuKGn/KMBzIVXnRumTtNPvBwRe8cL6B7wzMysPFiYGHUaQhXoH51WjN
BRWgQPsGSeupExJtVxU3nQbQbHMyAKMZtTzQTCUVSY7FRrALOhsyfsnGzASscWb4Haob1L3rs5v2
ya5+CvZlW1S/rqRtloH2igIKYp3nXkE3BcPzA58A41shnf4BFW0sQ+VTl0DlVffDFZ3tJQmVe/GI
kj6V1kew60oUGYvP5vr9sG5LxgPGdZG3DZGhqItQy6pRx3WVraZ4rd1hIXpx/tnyM2hIvWnTd6Ai
YZmwP3rwNxQqC/7qgfKkDR30uSjF3q6Fb4OvU9x+Rgx6y/Si9zSCZUUTcBNTGwhYhM3r/7m2xgtf
a9LsoFqQTpA/M+xTVyS4dxTjcNhVWEv5O8fQA0iGQVMwW6OLXWj5JonLhryvlQj7Nv7/bCnyWFWY
Y+y4qcDTNa7XaOouZ0O+HbsOFoPw4s8wYW4xXVqF3lD/qOLebIvWC2Pg/7t6+PpKDJys/BsEIwhp
OF4SCM31XRyxrUUqnZlfIEjw+XqmH5purg+yJsDBRgEtoIY64p/yeeJhjS3cVNvPeEXiuVcI63w5
uzuW2WmO81AuIRKoA1oI2C4fV7VM5l8YiBGNyNRaVKF7MyLgDmCpWAKaA4TameZ3D5RWcvIUG1D/
9aKHQx9uiQL2CxLyz7AqgZvoRPrxLiavuXW9x7oPz0/dr5j2ZsRP7ZEuYOYvcgCEws2FWrASS18d
iYtLCtwniin8Ffye/bYr84/23ykwdAaNHfO2c4EOXywLai2YpBtmgmEZvY+8SGeiRZAQ5g+AHWQa
ud0zXu9RjJHXDDMwVED72lPgVLk7QO3NKSyOFgG64pVfoo0p7sYrmD4ksVzAiP6JI9CLOnNlx/7B
rvWEQyrkYrouQzXVe9fYPBsMJrCQQJA+OXgocYDGIAidEQXVgJjeaX7m/ahr0FmFzaUz6CAKpc7x
dRkWJQ9Nb3p1WZspOU2Or3d2Kg4A3A9fRcHGpFjjKBSPS97AB21V9d6gTbplIB+BtBbb7LqV/S+w
7HcwJbtOwhdr2GjfimTb6YR4YD46BIT7oQh/PRI2bF6AYTIIaNl35b2Kbw3PLU9bJ7SC4P6MubVI
DUqe/uzIujWkPBWSAJKoeZTt/6k2gTeVVU2Qsuki9F7xd1RJnjW+1EciefzZwzi6wD4K5WwfYoCg
RO77XNAHLwr+s6vrMS8Q3Y3Npul9+K/js6UoN+cvRyRoEpTK0v3H7PLM5fLZaySN+3UP8FvcOMuy
uJLN/KuGokIZa8l3iNmS+m+Snrcgdot0gDdPJ2tRTSEMYaCkTwmRezg7/ti6VSnKXKMwpqdbWYV7
KfxkRdNinOt+SIei6+4Lhj0aGqTddJiqn2Pmm3eaqCHJCYKKQd8rr9RRpQC2JkxuB9tBUw0mmaiv
zkTPYrPQosHFHT/K30HBJ7iujg1mPfYmveayDLk06ySnE/hfKEarFVl79PGf8PX+tNjKDv4hjwhk
ePVT1Kg7OkaiqryLanKwkA3xsqhmywBoxHUbDMpTcoqElvkRGZW3lGLjzDqy8SEKuLDj9AaUti8M
8Fd3fULqlT+N2sV0DPN29g3T8f02M6kSxMAmTGfEPicgDtTHmlrCsGm1/Lk107i0QZxLmDbRV7yf
IPpO6zomBbUi5/DBnp80BFPFl/S/hhxcYsL+Qu/RJI34dCt7rvNtSnG0JqOCWeuyyylkRMmw6Bpi
cd22T82Qn7Tk4rm0qST29nJuHfo1A6wP8ppkPG+Vs0u8qTkza18qpnxx28DPP7gjF71ADwAIgLJP
vXxLTM51io6kZWCLDoSOZByyLAQL1gCl9zu2tFeK45rdIHgZWB5RNaExscUg3xLcL7NLBWdLIVdP
FrxF+i0oILxSfyE0a1OHIXR8fYRJJBjaelFm9I0F/FByrg7ZS8WLSUurTO518mrdHYMDbVCJjjyz
+FATPrFDqKnV9BVU0/sh/n+L6GaUMOInF0hiqzMv0I9ePlHKwhx10BGgW2rmViXNrdHsaUIr+6v4
WnTh/L66ZurP6PyTxXOiR9hZUFDhfF0Dnt58wiSCgr48SjxDE+bH7ykLoxNHLLV7uAVLO1cRXMre
QEnmWhhCcr9W8roIP8CFYpBZGzU7pERIKXen8oGR/jzffM0QYBCqomeCuIE6lxxWsLh9lcnJMW8I
t1Gu6kiksrQG3+xcnv5EgcKI6Yy1fui7BWb8iC6Vd2W0AkRYE61RshDGJXqmECWYdWxFoTiuWlYz
hruzEoqBYtYjQFiy6iLgOF3LuT7ftnGUOV3EX/8Kcpv9AAI1MH+MsFzZZdFDrHDT/Xcsl5lUSqDR
efNkgzhUNKVkV2to0HK35sHt7m6SuwrEKfwcJIAckqdNcQG31fjC4OPyI6G0kU9APb1v0wEYumj0
8YH1vbD98pxTW92o6fMPKkJt3BPv1EjQflfDBHzCFc7vIOB1S0d7IT5MxbKkt+ugXCjkcJUriGMc
4amvNNQBNrAKWMAk9UwaQlDQ2AkQG4qfuUMkP4jengz133fRn7miwNsaG8UOzSY1jK94B9n9MGr1
FgihupEas8PuJuL8Qxf5MNgVBvSVsykRM0+lAkfaCyyMwjpfvPzIrIavS/lyjRxRPMM/OkI0a609
qD1hJH+oSisocWxzZqOL8ZRdMl7yAk0Z2FW7WW2cRF1VhY0XKB25zwotNTuZM5WCTFUUj/QS0ARr
dW96nTzIW2FvO2Z+cmYqD36/tylCLs1pRvWPBXOTTxTTQPi063eTtUSfOvk/D4p+nPgBMslJlfxB
sbrqP2G8WKo7H9yTvPmlyxSq4lHXQHx9y4ERUz746Mo1r7miClaONA7pCIDsFHP4emybsCSyP/LD
CNeOut8ngIG7vMZypCHBEA6evgH6P0XAXUEkeT8bP56P1Zm6XAS2QQ11sl3ke+O6tgYbo50ILBUy
mvmAueDVcrTnh0Wsf5TkMXr5j12+JIM8xdzAA/k2d7gCk61eMshCBsVfTHB5rRS5tu7IrhGPLO5Q
JavGVWcjGOB2E6XKDwz6Ft+qKf4sW820cKS3iUYPJyc0TowBSVWZfSd8exPw8jz5QwyMvsMjT4f+
rtjp8qB9Ho9zccx7psLJwQqxEY6cs2fekLw/FefNWLwA60eriPBMqZ821Gio2i/bgkSGU74O5zxS
ChPmDc2Z3bbFREl6qwE+0TQzMWAvqzIhXGWmgC2V7Fe02wmED/qvM9mVNCXv8/lRzrBthNW8WEpB
ORBktdECsYAgqAwDZRQ//4d9eVwcS32fbCIpCaXDrIoAvl6FMvnNp1x7B9YulI6XY8w0MdRHKd23
5gsveI8PHjcqX+wfbCym/zc+A4cS3jGjOPh7Ysq8U1GTDpy00JFbmCczadrz4rhuqg93mdyJr68r
IL30TEEMsouQOYlYXh6ubwZNQbtnYHJmICW5GdF0HMxcvk/AIiZsNTENk6vlxCyKou4KXfquC6m4
MsLw0jSg/r2yl49P+MA3E/9aWub1JRHHBK9nJGB9vQMzuwgTJyu44FknIGTQb1ODyBqFbcR57jaY
4ES+vu/6n4yjQ6Lp0dfz36xcarS4OvieKT6HQXWaim4vvUl/fQFdnpphZ4evLMnf7WqCXo2+tQay
86bWdu6IB6m+5EOG5r5WQxl3fCsR1bcdbOUQCqmzzb3aIHoiV2Od5SB7u9sefjd7aLs4hW5wAD+v
d7KjtImY/11vUaqCmsfz4+NucPLJ4+setJXEp9d/DIStHWt8IsTJLL9ZruX8DHAFblaLWN9Ekjwb
jhBshfrj7c1CBl1lTZzUB4av6G1NZRk8W0zIhDITc0f+0nANd1NiNzUgtdTQjP2kHEnak3tyCeqs
HKHfTJKTNVxaBsu5+k2mzrP3cyQMitgHF3lGVI9R4q0Sa/dVOlswXskbWRD/xWnOxz/HXRy7U8LA
5WIvv0ktmAk/rL3JXiL7MjU5Zvne4A2oLSKl0RiSDUFY91ou6C/2PxiZ0NVyTjV/nMSfncev7gzd
kgF378/uCoGF3k5FqpagF/4fynfxD4eOn+w0Zd0eJTq3d5hyDQaSXFkHbA6szAAEqJYeC9kcRqHv
cHal9d+iwx+frvPAYRQN4z0UzavTckUJ8TBDJKciS3N3qrnjGMRxp9C9oij7GWfq8IV+G/Fuu5Aa
xCBgoTWtNNRDLla9TYwHcCkpiCieJUj2GzTpuX3qshFJ45fo8wAUioYxVtYIQKkOUTQOpFC9TtjB
aU2s7XuuOvUJkbzW9PAqecmig49hZRpX3nmaFQhrK1aYwJc7z16tMSdWT7INhZtoQOGvvgQSEyVG
zbOenuUI/lAarBTynHTufM9ZWNOngg7OSpO/TZYv/PWOtitV94n3ba6pbc8drarjSgaWjm7eVQL3
hrTh0G1AIW0gMkX6zs/TL+Q/B4uZO489mj79JlpZgdDIKhbT7RjwpPNh/U77rIykc1aesqyu772m
izBomBkMBQSI7/To24+a1bz4WZTdjt2qbRnLfwkAqeZkjLPPwDIyMVwYV2RGEE4VrrnrJHK/QCjk
rsnVq3wnsAXt5wihJ3j6PIdH8x3PAVBHnesmJ+wECKP2IgwXyCExNC0xHETCfefMOJ55HVG2bY2y
8J9ybp7TQGNIkTZcOYKbm3Q4JN7LMYp2tu2glD6biLxCF1DijClPS8bCdjax69YxyPlztjmrwM3x
q74Am2fmcnGe7aj+K8Cvz5BdRwRAtrgktm6URglhVIeSYQXMxbZaefN5hM0sjx8nw9m0/jYQDfS2
sL3/FNdMyDwt8ftN/31Uco9r5IKhBg7XpsSbmHyv6pbVldQtIbCCtvM052O107AaSrfLopPXIpY1
C1KGrD7OoTR4vmXXAxf35c3AvalqThiDmu0ZRjOVsUhGQ/tVPcLpqohU3pEKMA6LtPAk9SuLFR2R
IsWCjYRr5IylcZE750MaJjMvt0bucJOba8fr22FmHjmbpoEjpRBD2TqE588oNPqX/9S/lDhEc4p+
TEePHLpF2UXUegP/CcKUmP9AfBWMv5kuuknHH8UfxKKTFD4oTD8oBvrxG16++6fw407o7sb1aXl4
hYOY/wyhkokwTCILD8X5uRY/uEDK3BGU3bPDuBf1YBUtyvG0IWRwB/NMWpmmWiZL7PABWE3JyrNX
JNl2By9aQvdgCTn3PxmmWyT0TpD/lQDsoLOX4sbu0xrbCdsDcQm+vd2q+5HTcBnz5wtpu/f2Fi5G
dprHxasTM/BPo78uiAtsl7YspsH4TWrhXGyscMHRieQy13lJe20appbtMpktONVvCDO/0jiTqI88
j6n/BHRA6yxQjyvOERaB5xO99vQO4tAnpAaHd5aTWeN9Ewt2260pKVMVCyhEiOaXorbEl1UnbOZ7
h/vYSKS0Q7Ovaywgq4/JLAblMp4amxAX3dpeoRq0/1NlpySMmcU5fFNQgmZcOOfG1g26b4LSgUWS
095v+jB/blfzRoRNIAzvjs757xatXk0OOYTTz5XLMblEHEALwxjv5PCa+WncShPDLfMAP1IBzBJQ
T32Y8FT5OMOBSYQMmz3ECyz1/NKVQ1zEvbUCQytDBFz5voXY4ExuHh3BpLpEAkoK8ioMRyxvZvvT
kE09uiaOSC39Ba5klrHC4BzreiS5UZ2Yj302YsmUPnSzGlE7jqrUedkgWL+AsTI4f/wPAPYifRL3
2DwA+u4TVInWzr8PpmfdoRvkb33ulo+KwLH2dpmgPkH/YPL4e+Wom/qKDasdAaephn+EjyVLiiwh
xcY4+wcsYHx1etIK6eJjduQnHnl61M61l0lIA9oQWZf1HPirIlbxZOthW6FrfYBISSimnFk6P6Xt
p8/4U5TIhtZdTBsWSGZ9S941FLcWm4r2M3tg/yVh/LNT2yjiuT+GSrmfJz0QF0yt2qr286kVqyVj
SwSxd/CdIdQCRcV+WlSirwnAQOng6vWpiLO7s/2KfPk3+wQ/mf3LyeDC7rQsS7aGW9tpPcQP4V9U
1FQ3ciXkVdXj5XhR48e9jr8TvA7Tc4+cabqdKQ12oWxCtcZFPuA/nEdOOPb/TKD56ALQZqBd5jpS
2PtFfGeqxx3B/yCDr0nGTd1niyQei4QZSHJRpopdqNkuBtBUBBaXUV4qyNuHCt5Gs0PWqueEJDyN
9YixImKxm8JPiTJ2yU1Mc4ulnUsfXA51f6nsEGoc2itA4aak9ksEw42OqX1L/xEeQd9sqhkkZSzU
jGfoTfdsGADC3zgpsk0dRYV/G5noSt3vXT1adJTBmBUzppVC8qU1eo3vibJGdzY1pQvgV3tQo9Yu
UeUEgMIDvcrFmbdVeNW7kpzdaqNUmxcNh3PHGxK7D8fXtC0UUBAVn+HeU8RK4VHK6vBdrLxxc5BQ
TJIAXfEqYryY5B3fzHWtWmXukioF/gbdy6OvRV6k0tOWWjIU/aqmv5HCOVlcg8r+7+zBh+F8dFXT
bzb7owLOcLuNNEkCBmMGOxWPrSKqozBQcuNwh6r48vFK+IET2Tv7osW0YeOWeHpuJtw1KLR8DWp/
7QLn72/cdPMVZyIMHO5a+UsG3wUwv+8iyWya947M5ijcJbM4JPB6/f4fhz8gJCvevtOqzq9680dr
hYk5Wkz/zdhIGXAEpVnsTdFCPGQQ9dkhPeJfj+tt8RGzkE43gFNn6wbk1KHMazcBLoczK/HIo/Bi
4/FczkEj9Mh94X9md92Q9otLiJrMiMazzWScJfpW8EOFoMvBvfAlUDVY9nAEt4ZVjuMEQvNrsRa/
2oO/sBUVFMcPluPRNS8o+mgqDC6qIDzG7/zOIq22jepDCDCkHO0I2/BwtukkyD/ONKcEMGwpqx+p
+ymLJehJC+7u1rRN+D9wurPWNKZrRpSbFgpJfkHyyEDDHzCGfmeD6jREKjaBRqHPZyFqvHXJchgn
yZ0ORxkDGx6q9bIrADSWhokfl9a3qD7tO8v4MKzzv53c465WssxgZqcyiDPL1giZzdPfdgfbeYge
EPUgS4smsAkySe8rykIEVJp/mdpHZ8asw9jtCRhKn//YSNNae0mXFk+bWYeQXRTLYPUxnC4vAwsM
YvcjT6GEfcwaojTYHAzi17XeIFqfgLtmid6mxCZF4mQ7RGqzSMauKFjoqzN0xpSCYJkbWxJsOIdQ
Pxw9O/ntwSw3Fq7OlRxr95densSKC4bIPA+RB/yqRsl54ihhJJqRSOqhX9C5UpwiZKCBJeyF7y2F
4txpXOrY8CLqKjAWu12FJtAzfOv1sSo3KXf6PmkEuTetqJHAk/oclkNWWRarFWTPAxbjsEmJfjkN
0oPFsynCBIXJka9IpIN0iiqqhYKddBK4vtYyETdAOqkiEdA9PoJFA2HQQhMS9g09VM5jtJHLPDTP
It6qLutIoie4b7mubKLavq2e6WHphcmgSlc1eKHkSHhW0DvUpK+ruKq2S9DlpEsss7k0bWy4rEsa
vhO9tpmJ4H4UNFCbQ6+z1brS28vcaZtSczTdicvL1pl/p9fQjr9Sh40ObuwCvxWCXqLI8fwo16xT
LoiUyIIHJBl/WJddpVtsqMAo621tb8RRJFbS1TAyAiJCNgM8sEh1Vw3dh5mvTlyITToCX8sEM4EX
S4IwJaM6PdXSpvppdniiLyaMXwWAYHFMs3+etaZH395YOVmq1577JWHQ9XZZ7DMMJ6EMUm2oRbVF
GbQ+Rj2j49JnWjjemAU83wVARJ5gymF73GycnBix/E18+pwnU5pAJM/4ya4pxLwk58ou7liHJE+Q
6B+L42fn5Tyy6RuftDrh1Odhev9dzI/JZ3KgCFoEiy3IfdsQs3GT5ChSN6UgeNj0vIsSDdWkF2FX
1zdUvER9n0KET1B2F3F85hT+Jj+GSyUjY09pdGD8XPmn9oHyXU7Ev0glsKDOA09G/Q+tQUjP1N6z
BGqn2fWluycEGRWjJMDU+OPseGjDGEqQHkjnMQq2EwdFjSElFBQ2MIFdSufjOKHEKweYqvKR3HrS
2SjYm9fprDcdQBTO4XYBcfynhwNPBkUwSKRiQwTaKb0T41IT0ygODl6eBI3VhsmMAa5lvEx7+Xsx
NkzjS5IOHFq/zkm/1QV/aeGz2pYVzNsUhtd9BfqUfQHnFc8hQ1wc6sXgj9WcxYiMpq1x38BcGR+w
hxpQFtrxcFedZTpelCrkN7GH29spaZUMHvMoOKbkCgjqT7a+EHIEkLxCBydtSTS6D/1i8tmKMQ3v
C6V5+f8Qon74E0uiREkjo4BnvRoIf+IdY4pGTogdbro17gXMVA0Mn4l8YPLP2n98vlRQRoACAjXr
q+yzWW4AqI25oQ7LGSQeSIJ+7Y1tseavBDmM9gGqfYBNImDD55ioqXuPqBJmXtfPR3dIcbljgBAO
D7aN1mOMhX4xsU6jqtJT+utkPR8qeO31QY+1OegCaZM2uJuxAzvZZogvZZvElsql3Gvjs2FziWbU
pxImZYB6qgytwHXjoquNggyJhKViQ1RFzJ/jcrDzpvxpw1hz99FZjjhRfrMS6MqEbh6/pho3mXqx
7w5Vv60kKJMsaKaSLudKfyEndXXA+4xS2kEjH6n5IAYYvTiWXUVEUHPygJ1l5N1f7K8+B/c2hx1R
A7MHZL/UnJvssTEjyxN0UT6pcvhaCKfs7xye8V2VnTmksZg+5KXyUM+ArfF0eaxhYdeMMEgcIEFo
wQ/kIS/l7MkEKgyM6kdHUgXOnSU41f1sIKzIX+F0jZWB4JaRN/mUdPBKZqG5NEAMBEiPaH/Hy7pi
N2sj74qy+GOqnu6mU7DnS+yJZoLkUYuKUe5rCGFt9wTNrSy0MrHcTFj4SvsgyMLVS1razeRu3maS
/nbI0syFRr3zt2QB1SknPD/QjvCkXxzGyW+UOHxc1xqQpMSaCto5r4+Kh3bMCoBjFeGaqWo+IT4S
qiefSDo350a8e/HtUenaO0ws9JvML88wdxAAjH3jHwj4lOULDFX4B8Ucqn8kRy6oIBnwycMBTtHf
TjF54jsIWBf980PLdJvBe8dGgGDsKsyG1YHGfAs81fvlzlSztc5+BIG9V+25BOUIg4wJwjmlrB3D
HYz017QhdPVc4Qtpn1xofTZaM+8rN2LGOoC93tCpoNKOmwMq49BoXm74XEYlIJKExqs8IXFwYPKI
i3sNQniBG6kOsnvHg5DmmM/M3WkgT7b9w0YFT/XV6y8YpwKgBYqRJc3xo/Gpl/TOt9y7RCy2yoR5
b9HVpUrYpAVoJuyKkcY2aUWqhE8fEQuiTXIlqmodL5uku9DOvYXo/0Fq8ZOc7r7eeZ4ptg9AXmn8
MWLffEuyYjYiLbXc3Hem6zy5YnmZoBCvxboGyF6t6yTnDb69WhWBHKOwtfZ/UabTto3g/HZgv3I9
reZ5wNOIlu5LFp6JG1H61am0Hhq2nLscSh1R06wuwGzMQmC1PlUaO2YJNbOUaN3APLE9ch35eMlt
LmY6F8XF004NRaPsAfpnImNjIRjdDzATpZQJUhJyryu1LZFUFWRHmxCmQ8Cb6AqHEv33REr0vaiJ
LLv4dlbpobBwHle/Jm3BNIqSBDXBlaEcW0zhNn2YRF2vELg3eXEWA+zbBh9povHOo+PEs+bL5f9K
S+qK+5gzH2krJaOzd3jEpt0jGXV77TY70x02TVG9ChIlpaNTjtFraba3QeYNaYnZYjOQehtWNK5r
nAKV8kWPbmNljmdDzFZndP8BoJb8RsdYiRutsc3ISy55pU8dkvlT3LlL1D9Mck6FLDPYxn+8vv/n
s0dZx2JK1XaNJyHGr4tLTHica4j8sk6duLUkf6xzbky7kxTOb2njYriQlK4c+bTChVp2mkqTYC16
2aEvDgkKcvxQaeC7+ezxIaYh10yhU/GfxtbHlwThbBH+hwMtaJ3njsFMSM1LJs6TyG4OT5nZ7aTD
YnDg/IeSSkmF8V+kRVkKpvs+DpMjpln7WEtSyhLZLSCt4bKF5ssfN3hdNLsqdevgpnmdER3mkgFs
Pfi1up+bs+w7FqTVnthXYyMPJwbMAmwTiBV1IhJVKsniw8PTLAVW4tJrBzQTeJvvx1Ik6UXFqTKx
rL9xXeWDDEzlqsIDB0EtaLHTeZ7VzJiGuoKciw4v+6UhHwEV7ykpiR68C+agHIZjcO3Tjhe/h4ps
nDz0KVHAdayQ5MMaJ1ZVxl7feZoRaEW1rC9TtbuS3+t/4RBhO6j++iJjvba/TAd2z/pxfpRKFhSc
y1CyT2BxEZ9JqjrZEgy7VQ1M0y7/mAPp9Fs+se11GYxBhHzeTBUwjklHKyTqgBQIkwQkNsKVLXrt
vsNKgSM68ivy6JDpAbcUDrR58C+9eCIIkWEJHns7bRtn36/TZo4Cr4261FUjiB2LByOlyQ5SUTEc
FQa8bH+i77fn8teqgBxD16qKUfIO/mLdIBcGNHkRqjT1/rxTMIMSpeq9xYUgQ0jo3sfzNIy4rMhq
BkLNou8HOBqMPEMHxaxPybZfEE/B1gNGZlIeHW0NmSiBxifY0dlr+T6cjSsG+T3EvjsirqSwv9/E
LhQrWPwZ+NXgKs5nallRQBkUS7++t6QzI/8zGttw7VJbU0dg37oVx4k8oAnxoWCBg5tisK2PnJy5
AbDmj76oc1mhQGk6cB10s5TRan2uw5eDXoiiSoaGqGPNAHmbTBBqFmjfy5FEUPbPQCXtRCimP+e/
MwBm2WNYF7k+PfMaK/fELR6abziwGN7UTux+IRBNJAnmBxMIphHnBhCdUHNcEBO8BDQqjVgrJ7e4
zAjQ9Xw27cxnya+SFhv+Ompfhqln4fl01rQ8d8+oxudJFKZ3kIbfF2+2uNSPcUSH3WU0WZGfYEd6
YFxUk9uGrteqc1jr8cItSW+kQL1Sj1eH/SBwZcJohGeZ23DUjt6yHXqE1SpvmqMCxAhi0rfTlZkq
oag+KCU7ToDHlePwV7zdTKDwkoD7NegwkPHBt2eDSwvoK6Y0YogyCjoOetQwjeMfinYRtBDCz402
qXCDNKPyS1/UxLlxHMVAjuSme+9QXi+mHNaPaX0CZ5/rayvO6gYJrGAP4udQFiilcpY7ZhF7q/bd
fRPv9jNmPk+M2h5GcVRKjTKimOU+7j44hBdv2YTH10wXlE/e5IUz4/7IM1gTfsPGVtLQ5r8rXOSN
bjokEaMjj5wOzVb0DBm5qdIEQUGDf9ovR5pH4T5JS9rjaNd0wkuMUZDpCI3ZhxO3tV29cEdA6FxY
wLu5enoJ2feudO6ePW0drgpttdadDgTWqcmifSN5NpS2vJzVmVy/rn2txrvyVxAyQrh2W2b2oUGY
Yo2u3kZbWhoAujf3QItgTCIh5asXPWyfjFQZ6dBOKbsp6Mr/QTQm2q5FDqL1VVrHbuRO7Q4V7lwG
CTF28vkTtbbZhNkkaYzU6K+uNF+dx5NntdFeZ4wo9ltbCMUcEKsSZMEWRWOcB3hVa0mF/oaBPhss
KfuZjbWJ93knJeeFfXWKfQbpRXTHDTvXOVt399OyrmPSpdUZYjQAkoKps/1GGcE6J5NAaTqdWtAP
FsyzUVWBjmOOZ9R+Ua0ukl0Sd9KA50BNy0lxuhRVd5g75bTSaDG20lGWIcdVpSVYBlFcfzqlYpL/
IFTXHlE9Bf1Q9EGs7zuQl6h/IMhVSa2hW78lOWJeDPwqr6C8pYfZkEwo5Y0I5ii4AN0oGhJ3ZOhG
hqUoURguTHtvlFQl/As2Aqy+pAn87zXBQ4cux37SoHjeQXCXDOEFV+a5h4pD0YvjnBrWP+jriaMy
YUpAP5irdNBqFk7wprX8uJVb2lZ/VY7Sat5AY9G4pyLIpm6zkErSQXeM+e1GXbeT8Rh/SHgewmSf
ylmvo9BDBr6wyuBFxCBANXsZiBsuXiiUTO5Am3+/kKrV3/ov3Xh7d3xqgVgrZQGvaHXSPFf46FXO
EoT/MFL4n309/IXjD9O49TFi6OogkXTAVmaDci1XYIkvCyuxWt9vSrc0k+uc4n4aX6Jyyuj6MoZV
vLlwZUs1NY7KmNLy4LWtKZYkWHhZMU39VMPokBBDPKvMf+E5BYjOuQ1X4ChsOcLjkvhFbnZjlFdX
YS3CamE+oz2gB7nFnrZC8/dH+a7LMHjFa8uHA6Q+oV2r5vN9/2z0q6SgNIaCIGcLK2yJsOGAxE3U
+qlfanSsrgF2iahD35zGr857vvOg3tupY1V4mClfbHcgAR/kExPfkrr6GJ2MNIkIONaAp67kpRTM
4OJxiiQ4muSvrq1D5KXd3JN2uVNIXy8XVmcovAeFVLA8d7Yh2Rif1vEqYTf7UNlvvKBGuvq5Ga3V
KLYyhBpgHE0bGRjZibco/QHns/zPfC3xNskIQO/+8h3J9jYBNUO/2nrFGpdPTqPHtXpEGyYQW0FV
ieOzXa8hSODuZKt1zRMBZIg9q2bdBXD4G87AqHV79PlSx+vkCf7RlEE7ins93+/v3VNzWPr+nW8N
eYnsEtc8uGe5g3V6lAzmkDcnc0iud6nodKhrBAo8SFjXolxY8yEjG+PMScgRvogw57LpigUp5nkB
XgMs8K8DWCnRqYqDVlF06R5ZYqNnLSsLCA68SJGl8FqfihgbuWag0Jxkhdk7YlaxQ24OtloMuDad
JBHKWHH0RPyh13466gW3hL+Ob4f4VkPxg9RzGlffMn1oJwbAgGvweCI153eJzhzl2sFMefVR9z53
xLfWk53VpR+mli6SuK2rYey9dtucMIn6H22cSJXYc0FdPja9VJZNI62D4wz1PROmIQYx3avZyWvk
k9J98FPo0y2czwskzLq2d7Iy9VufDulNGhaWR88k60BzkV9rQLhI0GFxx6os1yNHeSxdJC5jcCCo
Mk3tUBh/x0wSdSx4xSN+IRQ62LsZE8dBVYs1Xa+Xzc4sT/51F+ga7T/JQAZO5J2Das7ogYK9Tz0b
0hyoReZE8p1tdGnVbEXe6+n81QlR0v7qDBElGZZziVzphlmMBRB/31fpzu9RbVoi45XALnn6MJRf
nDhfx6qhrXdyZsP8wddzd3LH7jsnFDBmFddUOAZPuxeqbyqyHrXa8MYgej94fk6FuOMQovyng8ao
Fr0+YelpIVt9XcUsFQMBwOTbAm1EWMGw1xZtjoYtT9u9WW9xs1phPeH3CLCC/Kt4wnmFMjEdR3pQ
eo42JvZvl3vgBYFMxXHiGtWV7R72f60TIesUuIRgJ8AiJlQ33WV2X+RmKwwRxmh4eWIU5KqvyjXo
XUmYeljUIwFhcgv+07mA6wVWQzCsqb78JsbySQRkMSk6ZdK9LwjSYocUogUnbDLBIRTf/bzr3KAu
oI2GRS6pGARwkos91AOCQYCDDA8ys3ttl4vEIaD2Su0EuAATbZ76dYCQVQ0bcDVGyV+x/4/xdJFs
g4lm9P31fPbXWts56qyrmQeAQIRH2TP2PoBsGOY0yJr2NMaGfnxibbwv/WHyzwSKV10V3QUt6E84
qdXRi1SXJjOSsEFqSthLomvJZBAal5gvfWg4F5PmD/Pk7fMszOTtT3PW349rbBR86WUGJczRWOnK
6MzuTz/GtlVoLD6F9rJvs8wQhFEYSZ6jztdW1JQtCq1H76Ozq24hEMtTkgYmuPhOBAbUjNR+JBRb
jh4iOpyP2PL4d9RazFim4tmw2Jx2llvyDeF8TmPWj3dMpJ/dObNPxgu2NbPXhz31Uildy5nWc2W1
zv3ZN0nVLBS1gwb5mp6us+puJtGTb3aMrtKI4Q3FR4XzLdVF3y7lUghsISqO09hcppRrH3SabY97
8iX3EBDRrBLu8HbHoDl6fed2wOtDveYpfhiu9YJU9sbPF3plpwf1CI0CKga3ATzX/l89Rk9qVjlA
VpHZImI1QVWw1ljRGzwDmaH4UZm8u1KrgYz1sFYPp3SFEkfJND+0EMtbekb0YYZ05gwmBOK47XES
0fys2dwihVDl7Sm3ziyqogIDu9D5daYE3aM57zRX6Y7eG1+s4y4CoKPMENM5Ma1Bp1o2u6yEVJqM
LuBCwtuJ2NKof0KZQK73HIcUb8ctjv7AsrWy4xsjsN5zwSYwMfzFyInb8G+XBL7NSYgCr1EMOe2t
dbFB0wYN0CZ7TIZgif36GNX4Ibj+YGqeXFBzR6yHarV2LRKdiui7dL7HZjcOga+wpl5peZOn4Jnn
8o7bgAA5Blhjm5frdO9lWhTMjOdnLmA6H9rLOP4xT9ve/ZARl9V+HERm6nKHZ7Qi3LFnJlvGdqmv
WVRFCs1q6ZW8pbkH4oicMDU05PRbaovctCa1sDza8Zl6Q+k9nSOEbS/byGRdki14Iw/6trWIFtTG
qr8KAMyz/PN08D9SamEpv/sMaVT8g91B1bBtW33sWF1nWMsp3evIIKqyzRWOf+H8tynvWfrwadNP
26MOad0/HQOAugO7YQmK2KY+ZqOhrv4gDl29jTQyPYduUBkEZpQNVEM3M4Uv1WlnwJyZjWDr0o2/
G3DVhJI7h4l7DMKH62dFQsG9hTOUP3oBBrK7DsU6YEoTLrVa+rRL5gPUiY6TVsKILl9K06PqSkZs
NCC+PcdI1oz5CKK3nMa5v+PMzmUssiCd7FQxDyI+h9MO5khzOh2+R1+AHeXZ5+bK3whceOoJJyk6
GSPib3lNKiWfFngU+TK6L772lyJfh6qW9yQixnzIPJxtbwDj4ZObtktRhCoBfL+Li8EH/rsU9H87
kopvYSeFVDyGf5HBNPC7tTleA3VInrkfvSyc/y1SW5PKgapl5sUb0MKyNQ9k2sFxpIcU5Vi5xL/Z
+YMyhTvFMm2aMDAoiwm/C1ydDqb8m+afzYho0OlFcbzU/+egmW8jOBqG8f/dHy4fAsgJa8hLTbII
xHsfjxNEvQYFipODzqcDuO5aMTGeH4lo6E/NERuEwgO+3HEz898758LJS1KHOAUPxReT4XV0sjj4
ruje76sgkDJqEnVJ9pyot1ooX3v3z5SNjvGmfbHOW3FPslnDSbhxwXQaJLuek6CsgfIVNyiPxLRa
XRTK7izCLAvxZMLmvCrEAW0R4HeN67tSPV/aB2CSXTaiUse+xaDzFq1qONVzt9ML8qI15j/gi7Vn
zgyjesSog08TJyKjE2AG7K3rUptVgBqmwCpOaNCXSxYyFuP3cPSkn73BqRftAzNBECcWj9z61dPL
i3GfeIrCcqqxNAXgsWb/969q6JO/92kOk6nCCcviXtml8udpOwnRyrkz9uHPunV7HexG4QgCWkYQ
/zGtmKDlklrbJLDHr6G+uM41Ic2OYG4cnVRZIDKYT5SF+4uCAw+mi5AHKs4yBb9aa1JmT7Qr/o41
rsg1DYNqEVTMWg8n6q/+tZLApFmvvZTBLbUf77xIC8dxGNBHVi1lbvlWqpeSycmEDQ29kwgZ/HtL
Tkqi8LIx2Lqmhy/rbRoaF+ypMGpAAntlp+AuV2iLRxtYx7RMKSYJ/GROd6WDAa39nxXbf73jiYJ8
fA8AslM6tYbigjsX9LZNKq11K3pV2Wr0GjZHR2s7aEVlNRwZlZDDfJPNWBX2UIqFAuY43Q6jzK/J
KoGYLCvGUbedKypALZNgmRn8wTOMnArSSVnA+UQU1wRkQ56mp1ZPGB2LaBoUpHteeVbn4W2CGvLP
i9507z2Do6n1OkhbXdHZyrBUgy883LdVZcysZvuY6FLhVddVh+lkAD5vzTUC5UgAK7gQfrKn2/q6
ql2Dgfh3Mw1kQP+UKkNufOQWJnpnVbpdfnQmy6gDOc8FoBWOWq/75Pcnm4NkiGG5WJ3LnOxla8Du
ORF4SIma8lGNhm5+hCLxJ2ZrdBVUo+lmPU+hcdMm+M+grM5nHLHXgzxBbF7b11TsxwS3cmtrPu4E
hOQRnKATfDah37ILd2We+KnWUSHf3wwih7k2LWnjj2SOL9BZpcjisxO5q4I0kYr9hYY8K63IP1nv
vknKIP/3mBNg+bM8orNoyrw/KpHzYkYZDCQOL0BnpLdTRHwQW4HUNuMbWQ5munNHteMU5/THHCcN
T3KdtRxlhZYWYiDZ4MCp94aTe7SLSc4u7css9fCnxKIFegW1dLpKQvXh7zJrGidb1dpaSGupBnAl
a8KDR/dhrOYIWKB6XyunwxeFZuEHY2ue9LJmAyJ45Ap5/j8nAna3Oxqwunq4aTUofWh41LD9oXqp
wjynbB2GW6HkA0L6f3cUdLK3ZA+a/Gcj8obpQpqZAoqw+e8kzdMdQBs/xrbN6LzTkjR9J6r4SPrM
VTg1iFIEagff06BeFaFEGy4yb1pChC+JlzS9Npk90lcIjW6CRT1DRJR60zI2oxvLedoS7NC/cSYR
E3DKJzZg7DcLHonwylqLSjRsLg5niHTL+jqAxSAhJpzuGel/NHqZiWYLfyj0FNUABKU5NHUaizq/
OKl3g0ck1SdtiwvLWeVumt27+w8QsgPNxnPB2cjJ+QSgMuxs+Ax9GlK2ynJ6F092qBTbdHtqoHGN
cBLDCqT6qJJjrCRqi7/osbjXovMpj0A47sPhEMySvGa6wpEFTkrCKa9i3PuZmBZwcHzwdJAUD+YG
qFkWGcSOVGG9CUBNu2vZtLHS1cZHddbFnl2iznI/8SGb9TIwMGU5c+0rp1pjEs04aQ9O5DID2He4
aKCO7SY0ddt2g8fDcBaPzdJGbJQrM6Av0db0CGRJDE/77ljtr4wxoXFqXJbhAGIgl2u6uOC5mcDD
sR6107ADhjpUL6sF1JVtkUn5FN5zw7RJA+Z9G7NT9d9bJ856Stx5503ASmnBK+xgdJsbJE8bsSy2
lmKkz3h4/aZjzCa69St1BSdXhdIBH2EC+bcvEPqCpWLA2JxZsKxbG21G1rvwTuXMY5LZcKx5Yv/w
76b32ALkK3VruspZKMXbwU8toCvyNg3IPT6iI00kJkjfXJDvdx8roF9n4uXh28CvgrOjnRSa2jyf
khaPdCHM8s+DuEEeW1PTv/i0Rh8NqocT0zfk7m2JR+2pvljUyniSjtJzf48v+72AVPE07OTG4HiD
VhvKKgje7/iKk6M4DexM04ZU5TAwf1RHkOuJ4yNTTn7fLYkOdqzVOty5SjIe+PmIeIzdMhNhjntV
b/1ZVWOqYHHZvMlfD49CYKDf6dEID6hMhmTi8p8K7mXt81B11amspo9vvcjZOjP1YoZzvxikbZZP
8Fe0ilsVVzS7yJ6j5j8+0umGs2+Rt/5f1cYrb2Zxvhvh2VBd9MhyyzYVd+68/pVZTPp4TkLnnvDZ
9fT1K3PGPpSjMn+6DyDmwg900apEYY5FBZr1IVb4Sdvyywi6Veswx+b9UWHrCnVK3CjLWyyfk/Bk
KOGapAGMIsRkJ/cnTXZhq5bIaFoQTHi7tEz24+Bi+cDsNngZjmcl8pKgbfxFAQCsIab4g4i65pyo
O+IJ+UpQGAxCMbTFfj01seLFWYDqC7WePhs6ptK+ui1qqU6mViCqgtyNxVVtnfUnDfC/PILmNkLk
vkKQBQ9i0gmKSrCBK+PfLCm78gYvphApXVnxBvxbTlfbO9R60LUEtl4heseV2kz9PSD30/y7xLXT
sSIiNo/H+bqsXPi+p+iu2BkX9KcKYr07FcQzGg+BnGgB3z8gbw6NlndcFh0jQiEKuvJE7NS2+DW2
V7lzMRg+gw7IX5K96ljHOUcOEoLa49XnzxoHmM9i6b5hnh4lUl7+JliRIG5t6tqzb7h5GojGd9Jf
JK5lH1ShGxEFQ8F+0PG06NQDu3WuycY51R14/C2TSFPQkCrG6iIzMNkFpNOakYbNHLDVSDDkAul4
NNDosCTZhaVIZeHdHI6A41uwWP5q3C/L2VT5cG698PTwCzK1LZOw0y71OyHlHbPn2XtcVYb/UXBM
4zpMDi44AljbGHBlHPGlbupi9sTYVC9PMNMk1N4iSjhDxGzE10A1ZSgezvgud3mvwx3OKVzcZDPl
ZeS5lUPV8nv2oQwedcHmFlqU4muB6IjHG/J6dfjJiQry7qRLq5SKjF0EAaFMaIk25Y5tsdeeT5vo
XYsWjxf6ad4PwJyt8hUgWtuDpUr64vgiHENn5aryPt/pt0Zg/sVSeqk8IgPAGI6LiwWshzUD+F+X
m7npo0Wa45mDFQ1cG/Fd0jMJFWcGSHJF/1ssCKAphk8v3/iw03xE0b0K6FGi6hYy2nWbCL2cOyWM
JgUwdCpi73Nhv3MrWPPS5T34EUF4/H4/M1M2x6FQSrDemto1GmEf2A3zV/VXB8KfOWJfCqys84zp
NXsJrPNeWOa9p9jMtPiF743x2KGqT53EQtawu86H14m9hZwkGKfH6fOM9HGXt3s9Ypi7GyitJR15
FY8cLLZxP8ciJVmf/Q+cK/t1oK7yfQgdYiLyAaFiyhssk4zON/d7nvYuCJUj3AvbOeehPVf/XZ1r
8ZPENbY157KiVQXac0kz8p6Ynj6I1hMsf3YbcKgPtPIIW6sQqouwHTPkuaubdCiZFYQvB0muY+/a
xRXgYGCNVsnHdUzB8opkJiHGRuViOir93VrEqWPkRzmFwUa9FvkLUd/GQMZs7Z2oidzaDPq/dvUC
Gp3kQsLBBYZC+6+7jkUj73tFMtYQXRY0RJ8iNgmWkfW1W3n+j0CeiEil3VLpS3LloGdLaeq60lu9
VsperFdMqLM1VK6Ij/7qTw1Uwqf8XxKy2hQXPMKaLMwklGC1zfiL6912X6rSV/dw0283tB8MTMyL
3HFDUOlwx/nMS0d1J3wEs+ER9ZOXxgd8DcsShby6uSSTYNUtmnZY23LUPjfYU/DUeKtEzoFudZtW
ALPuzA4P+4hkEi6u+3ClI8bFYrNT1URaj3kncfa7GUWm7PdZ9ywfEODJgwePMrNp5QX+K3isCWo+
cfF1ZMm7FBcTJ+we8cx9lERSqVhlCgfXD7eHz4lZ7HaleJGg2sIfPB6PkXRPLQ8BikLSUmGAe2rD
ecdcL5Mgl6BvrBbvMbVKTxFqaSQr3fdRywnr4hUK7IQ9ZGJRe9Z8YK76Wi+BG+lzQHCJpHE4rOep
wUJZ+sYojGdSBT7LWkyQ0LbGorDiuO6V4I49PBFcTJ3cpJjGBmmJjGFpwgpx3nsC4m85UhNrjeaU
yMmtmfdZGMeLQs85Z9Jlebmre1ODh2MKLg+me+2B3+BqxpwvtqCm51SIkRVMA+/882i5IDn6TeP7
ZTknyijTOl426G5w6MFSugnFvjLTEYP9uWDMmbpOgqyPYSOW+ZBldvjQiDzfMLetYGV6wmXFAt9N
Aw6WSICrdfMllJ1WxaKb+izOk8JKwe8Md2DWKn12LDzkq4s7fmqbNGurHeFrNRgb3w/51ouXlDgV
PnywkqmguekBUspDepwX3BvMOWuXRjww2YcX4Uro2UU2bcPSdWkApX5IhhtnStsRyjo1ljJKio6B
DY7M6vuUZmFzRGaRx+jqiIJ5qX5/knEYi6qllZ8/svQdMiEFMWclrJjzTUan9MED2tBxyOHaWGtA
Ps+38otE5Az4GDo9o3nN2IeACTXItbySepvW8veMuzkesOB4kagdkdSyuZBChIXFie2bRmRanX3G
EN5u9nn0OQq9SzdIy55394+O+FKbEh9wFcKUAkd2boQWtJRcKIMwy450d4/mgfLcDUR6KNJHCvte
iC51aV9vEn8bC+aDSBGBZ7KqyOwB08+QImh6HYsaast07QH30oSYSoCfcQpZIjXxX/G+uD2dB6So
Zd63lQPV1AzTyerRZEMjtvkl3FRBwOxgBFIoz4BBmmEm2RN/Rn6Cs2WSQJl7etNV7q/a4x5apy8a
Zs24bmVuPrE1jnF7qKVWpz35tjYSQ7YMbWr2COUk2XkMt9ZXTtOrTbaYDJcEgezxHuKPsFV39u87
2s0xFagcMn175NqXbdp8PDAp1VFntMbkgHufJ1khleWcL5oXAIwxg2zwCIE0s8q5FjvVj7PWP9vH
1jlzp5RUUtm3Q3uda5N/6NU3zOG/QQW1JCJs5AdxlMCYEHHxQ1OsHg7kBziZXBkD4sqceaSwjZND
mBrPI7tZXdzh8PmK26Z+JEUcxl/dNhbTiu2gwNxx3kPYL3HDgcB6bD74eZu5C5mS7j8K4d0Ro385
dk9dcF/fr4atzRdvVIK4OOjV57sUos+1jAPQgfG98vWrHtX7vmDVLh/ZUP/N18dTtopv/jZwIBKJ
72lpVCAi7TzgfSXen8Bx3NpRCsdIkpixhkIesEFLZiXTQDqiDmC5WnCNIBbG3TvUr3BvSxCanj5a
/+zqe0MlfDt7LJpi5nleS7INc8CwdQqjGz1jj1SvXAY8dOa/1geDNEk8ELU89yTuIoKMtPa1Q08+
ewh2pi40prkFPV6WkGuykBH4UWZr9I9MI612Uoxt8NNhi2pBpwAbR2ApkuGMov6ti8iEmL1YwbbS
dT9rialiH9M/kMsTaqO7Tc+s/1V3wotulY5PnAI8oDhzGaG7aFsZiS8uUBdW6JeV+zuqR6LE1kph
3yl7jUSApARPKbYeoCjwqWZcPkvwlU1q1+oo0PrXXZSrrP1VZ3Qkzr0viJRthkdWJdTejhqFl9gj
1i/WAljlmkk5Y3bnYr+774ppvAE/pNjB9mDHMPA05z/kRQwxGV64+IhHMtoYH3U6RgfoQesS47Pb
WW5Kt2MYfH8xi/hSUAFsw+MAX7urCQI/yDuyn2yrlknbX9KcYzfkuv5AQRdzJaJszxAvL56T1SPD
uRnkds3XD43dq6wDWPyHsvw1TuBnKRK9fwwf2sstsyT0q9AHEwaSPdv9w/KMSnxsFO+Hw6h6vuLr
bDk23GgTRr99dd3ANyBWc283ubAPe4FTQRdiUuINe259NneijGY/FAyrNrnqTy5RsaGuR9T891/H
veDPqsfDqqcJJj3ZDHEDUxvogQ+XmlnhHNC0l5nZZPb2U8Ocaoe2wbWGwqTzqq5Oj6KRntW2/723
v1/CMlZWOn8sY0j7Olr4WUKFmVCYdzeR/wI1qOKv3yM2V+XBf/m/Vvh7ZpSQOQ61TLGJWxZ589p7
TXGz1nCOWkP0M+eY0SytNurLsHSePTpRd5t0rVbTXWZZJOwZrCg3XbKWwn+aNhRxwqyrOurwhMf6
DVW4rzIFLM1sXt55rE1Zhx/05LgOS2yLujFEarLHvJNw8GgAxEEfx0JjcXJ2GEJvpINIC32Y/Lpx
lGTefG9JqozVl3uDcm1A5YZE1z9PMMENfAZk3g1zRZVNTDrqLRDRlYMr/6gGDw8jLdslRBpWiyph
Sd6xTubNMVnm6rPYVSkYx3ftzkLNhu+nrFMUjpd+q5Rn/jbDpFF6q3iWFmjXkM9Mjz52V29F9pVi
ySKigC7iIwVhYmOmplziOHQbnRA22RNhhOYyRSjW1VtpWqc/pk9ijJtlQ29CuZtkxwMU1FPLJ2Mm
XuSceuO0GiwV6OErStfZYSO/9n7ofjUWuWehrRonSkHFBiQLzreUCQXT8O2B/KuJXY/DdVLpH5iE
jpWuESLIAHqlaOdU+sCbDivVSxYlgs0p9DZHz8UN3CXBTgU8eB2zP26RoJD01YBV7UkEf08Pjd8H
9cGGApmgwOATA4UTMfwTAie5bK+LFY/OlEXvvC5ZLPNhYZTtoyc0yzlICs4TFRO3y6qFF17vc4xU
+Y3fQ14jz4r6Ov8bKrw0SvvmmFEwI3eal2FMrWn/bU+HbaRKnC65PjOAY9yaa0/9iUaYCSNt817T
wdKzUTHUgK1A3lpjdIKMcJqX8qcz573i+X75lEl60HTFNShgE2iL627OUIEDc3daYeqg+EcZbLtt
CNe4srJ2YuZcqMq7MwNIxeNbkpuW5eZL4r4ZKJqk64OFitOQg4+O7OKl45esrlTlO5hmjsKsn41N
H5jJ8gFRrLkVo+/FPUh45aoBxF38DPN0gDGxKxrh+ENxgQCeWJ2iKgEqK1LhwyqgyWQWlKVFV1NG
bf9wU/035to=
`protect end_protected
