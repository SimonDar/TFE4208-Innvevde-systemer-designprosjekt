��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��·t����O�ihY�p6֑�1b!o9��ZA��q�Ħ��ȶsK�4��_M�s���H��`��c5e��"�X��#ƃ�pB4T��e�F��q�9��*�h�DM��L�%"��_*��&�AI�_cC�����7{�R�,_rB��_(E��jm*@��U�1������Po]���؝:l�qřː�*��4����s,����]`َ�_[8�!�$*3��e�@D`Њ4�k�l�4��&��w9w5�3u����$l�����sW�4C�9��U�[uSGj	���_+��ímL��_�g�D^�l�i������v֮��ق[|��B
��𼌟�ΰJ��2|�)an���Gb��p����ۣ]�<�#O4{��[��b5�Z���o�q]���W"Q��Gi��?�����.L�\ e�����|�v��� jw�$�����- ;آח5QK؁a��/ꓬ��P	��2�~PC�͇��UR W�'2��}���"�I�`�=�����S�5��0F'i�,�,j��7O��@	�F���.�Y�p҉e}h��W���@l$W&�)U�a`���/Q�д�L�ꊦ�5-��aD�/�%k���[��JEF��ϑko@�V}W(9݀��^����O^��F#�۸r�PTa�_�C��/�Ӡ�7�M/����ϙ��F�ڙX� �����b�{-3._�1'R�VF
+�L��,h�s�ԯ�0}o7Jӂ�<�*A�����9*�jw=l�����@�,qF���|�:.�6yŸֶ́�!�6���Mi���p��*�!ƌ:\|�u���W��XI�K/��F��t��#܀.�bq�Z2���ῌWH�V�E�5+�	+�������0x�Z��]a��&b�Eˆ�B�nYvgRA�E�`�T�ͤ��zUݜ��˓]*Qyryۢ*c.Y�qB�q8Y�@�F����U��
/u���p䚫YhQu��[&�����f�k�D%�}V��0R�[-@���2'�c"���_I*�-��嵨d=�x��k�چ:�q vJ��քou�\��M�ޤo���X��$�xS�RƄh,��~��|�\��\,�mJ�bw'��+�~�������|΂�?��U���ݐMz�����@��:�_bI�Y�@��/5����G/$�|��a���M��LW�U��L���ŷ\�hRm�J�%�j̴��>^�h<5֛:LɆ�c?���+La�A�����[�H����'�� /k��~`F�����;~�a��E��ķW�7��KH��lK��������$�T+L�V�ُ�uZ���?��D�Sn�>���g�g$x:�*����S�l�k,�T�S�mt̾� ��W߉�W0�JR���ᑜ��LßNS��Ca�|z�g�&����x��9����Fِ�����D*�.���]0�#0:e����3;+�D������a��cڝ��n�2$�(�`Զ-Ö;N�7{<�̘ 	�{𗎃����3��O�u9L�ҴŦ��1w��E��v�6WYyd��p���m�z*Z���ғ,��O�Q���M���]8+M�p��krgڎؘ����Wa�t	J�5�B�V	V�6)�	S�E?1�B�G"Z�h�h��� T�q��a5�yS�9D����������a�m��~4H[�!6Y�5��#�3�@���/��=TK��.4Hw�WI����`7��~~,��-p���ϰ��`�[s+`�p��7���ཧ��.�Rz�ZK����]G��N敝�����N��z��[/�3��5�8[f�ϊ##�1����rҀK�G�%�6"Z��6���=!�]�tr뀌��e*��c#v ׳+���R��בYJ&m��G��<�7�$��EQ/}ˮ����*��`"�R�t��?���*3�9�6���{�`��1[��A�ąIt���L��(+tuΑi毚"��zI�����Q,Y���F����\o�:W��ʽ:�]W��cng�F�~V�lj8ͼ��Π���d�6��E��p0&�	[�^е��u��]�(��rY���4�T!�ij�8�z�$�0*��\�