��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~	U�_K�-����(�谝�of00�,�#ʵ�r�d���(��Ҙ�[�Ъ��ԯ�JIr�*��^��Lq��q�	 #ב�D>�gZTHiꣻ!'0hdU��*?l��B�Ei����Mw��D͇���4��|��HjߐE��C4�*�M��p�^U7S��.�tz%��wQ�c ��)����XQ;���ϥ�g�[���v!�t�i��y�9�T'-2HGd�)���^���;l����+��m� E!@Ӌ�[o�K�3�پ�Z�!-�US�q!
�������m�ME��$8����~����u��l�A)�/�ѧ�q���c�����oN�����̐��!B��^�m=�^6���p�v��js��V{Ss�;td�A���<��Y��#E�^��%	���~���i�%Kk��J ����B���=�0����`��]��\�׺xzwSwr�'o/���P6I��̉�-־��Ҵ�G1F��:p�d
�_�G�|A��VokrH�u�D=��7s( �g�n�z�@W	0������$�D�L1�uf�8��JL�s����-�LUP����֖��U�`a����S����RU��+�趻ce���I��ph�_F\�����I^bu�kWr�N� �T�;���᮴�D z�NND�m�FB�G�L
�I��V�&�o�ɴ�w�0t �>.�1e(CE���	B����w)����m"���֋�L�G�3�.�Bͣ�����@�=�X�+�*�괐�����s̞�>�ŷ!$���ٯ�c.f[Ž�g�䞰��y�
�D�}�h����>MpP�y�a�,yP	�
f�>ԭ�^ɤK�Y|�ZQ����>TB��[�p�=��_Q�����=Ms3�Ћ5����;��%axˇ���C�l:�ڬL��
��/䭅�(:�S��vb�q�r.{|_���<Xm�.g���ji��m�a�cms��d��^{�<�ZO�{O�D(�b�!C~�J��q0K	8�CE��q9���'Y&�n\�����D�'�z�0�y�~�N`�o~^[��}�0� ��]h���ϼd�����I����%Z����Y��ծ�4�L=p|��JH���N�ҢK#A3kCE\�zU��諓{X�v��g. n'ujs��&�w�ь���S�)��]�c�v���z��v�E9�F{��֪^�����.��ZP���e�(�G,C�UێFم�N�&�E?<����^�ѿ
Ij�}�Z�o�|���*�R �%���0�oZ8��կ�3���ӍF�q(������x= {W��;V���L�%@j"�"��<�=�Q	��b9�Y[J9	o6KQ��q����X <�mN{�!� n�Z�^��Y��l!������a�Mн�����W|%����Ԃ!���+�DYd*���[M��?U�r-�:�u�[T�����Н���
�^�@ ��%�F�ӎ)��+��+��	d8��cBT��`���
��Y�ל����G����!�vxr)�lި��P��'At�9��'�/�y:�ZpEA���\km�;�8 b��%�߿����`,9�O���m
��V�j���r���=�J��{�b8x�hQ��z #���<�>�1 ]�6�Cy��8u=~�&�`���_���������>�G1�Gkw��� 1��)$�{��8z'X��~n�I��ܽ]��=�d����!�4hQ��,N��x0g"t;Ӡ:���R�%[����-���C��0�P�?Qi�D��>�=���I�������z��<�+\�/�ǭ�_�(��p锡I��=��b@��IȺ����)�ܯ�b�[��T�/�9��-{��u��4��`�~AӁ1���f2G� ��)�6mR4j����K��A�b����v��@����o����),��#��B8��#�ǘC76}d��W2Z��H��$�4��XpF�{�C�>��+�M��m�f�7膸��o}$�� ��W�Yl�$�H��%���/"�G,��yG��bօD�ƭ�4�7S��v+�~i/\K�7���@[`��o:����]�¯�І0�����sHJn� ����1����1����Բ�����u�.�ɰ�v���e1Z��5��(r��� g~|����e� I]�(g���őV-�Nk��NB��ko�ր86K���m����!E���<�(7`����#���t�X;���逰b���;�X�p���/	H���ı�$�@��ImA�!���~m��Aw?�;k����0�W�=��AF<F��n�f嶺j���ֆM	��¾�T�[��~|XwMMu��1�>-�~�;�\e�J��A[����!����P~,��jW�<B>�zv^��<�8;�U��kH`�n
7�4'V�!�5��D�p�#Hv��*LD��^ݐ�����~0G��Y�n�w��鷼�AY���K^��Q٘E��4g�I���H�6z�my���U�D������&��:�s�(F+�!�j���Z�+.}"3�maV����|�ir7�K�4��3��M=a,u��f�ѣ�����])�. LA4w�nj' ���9�YZ\�"b�X�N���*�2����魘����Q�� �Z�G<e��`bh3�7F}Ku X��%5T���=�`���{��z3 y%��gjBQ
��0����$C~�ٚ�1�r���&�oʧ����o�u��Č:��|XN��-�Ӯ���(FFɶq��J�9���üu�p�Qw┦u����\��م��O�D�Б|���h�'��R�tT�g9f�9cD`�,$y�c��b�Xo�SeD֪m�=_DNO�"�@H�hɁ�^�;�kr��PP�Hq��6){S�L^PT/�
�LP/I��OsC�����ZY��e���=��`�"�w��I�uE��|���e�.�+�^q���:w=�����{�W܁�Qv��Z��w܌
|UI��p�����6�It�����H��y�'T?���)'n�^^��S�W��i�]ۊ3g�Bv=ф���1:]K&�Tߚϳ�r�h,�3����0ѫ�wu{iQ;����$����	�t@�?�����0!�}܄����������"�[���s�k��дOm�������MX����#��$ve�<�'"ۣ�/Ӱm�n�y1�+��i*�뼤���
׊��4�Hj����5}mZkū.�ª��>!�rvt�g��dhr�A���r�er���>��h��N�⁸���ؿ�b*���(ɕ��L���+=�V�ąn�N����ڟ���l��v��G�-SQ���'G`gl�!