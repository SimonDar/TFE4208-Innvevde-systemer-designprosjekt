-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
l0ZKGTr+RZq3/j3dXBSZJ8q3IQdbuoddjATbMo57dDhC0U7fU9BWzczEOFLmRtXLhwjhorqBSk2N
Ml6yYVdcAlNsi53UAufehbBdy3QeMDlGcfUnIixXYinSUyxwXj+AOG9w8atJXyDixcdMjSBjg1eO
yBDAdw6P5bt5A+vcBgsUnbguDghJ8wkVN5b3+k7OErOtVC71MT2IjTc6SLqZpWajuQdIKo3BS93u
OqvU5oSVdu6RRGNFZuhsSmaOYRG8MKZ+cr2v6Gr53SthN6NXvzPhiSNnoxgd9r00GTMArGBDzYla
PmzTElGab/W/Ne/khlY+43dsKVeWBGoajabIkw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
vLB2rlUq8+irNH4yvHhCgPiKwQkO0EXDyIMYEexuD4ou5zIzJR4htrpUOngwsZN9KkPJziQJD2TW
bYRi0VZv5hdJ10Op+nI7PH4pUtEguW79h1GTsCYe6DH0LedqFNpDEim8V1I19rUZuPCriHA8y44R
tSCuft4GvCxebgqLs/vTtJ88ZoF/v0Y0p/CnbeFDqN+r0JpKet5Jhk5r10iAFVnm8nzwtiAksGw1
y1IfgOyBld6i2REbk8+dq3R8AySfyDFxhvete1mrDdPT31fOJOcIVO6Pobu6ep4IuMdv/bIrEUme
tEuhUAnHiBUiRFSz3K9UPLMJQNbXvdVjIVhVytND9sRSePgAPtsbYc6QzcHwgbcN9nwl2WTR2VWA
3FfFvNr38jPVDdrZusWjPGYNSgAN/FwU85NbUHbeP5T+9plzbSrmlS1vID2xXbwbVulIzrTomdtL
BBR/gSWSe4FsZ6zUncaTg8XNPFZyCumGDjCGYJJFyJ8rqVh/0Lm0tf7L3IMQecoLRcP+GmU8Zh16
4LgkEayChQeDK8GEi9Wxx0/0ih7c+/9aAtyrCTRUUWqs9TQGAQkEk1fDfFXADDAtkwjeLPi9Db2D
bZP6w8N0v2mSgH6/vM/WM4/yLD2PMSoqt37fi4Ra6QYKW5+KVqLsIS4HPPIRxoHkFLfBohzMiW9y
rZwmZjn/n1GfAF60w02PxTSV/ji1gHwylEeghob/dSfNqkf9xt7eHvpoYkYcuNHNtE2vyed+s6e3
J6hB2bVFhoAqzfz5hYUsoUa1bY8AqkA3af9w2ap+gZ9DaiH6xd3HRytnvZ+NbuLxZC7r7xf3uoaL
l2hFvFqrHaiEpoiVQ3U2agJjNNmPUi4+xZUeW2WkxyGuKxYwUHfDgwdC/i/T0KIISIJQE/Vsphto
SgJlDKqX5rTF+fLrrF2Bv5bYjWnypKA9IKUGl7XEFPC7BjpF0TAfIWAOgFoWugRa5TpltF4eN7Jz
5AmoNscWsJ6LrU9NoOLFgMGFHlNOirCpr4qCb9NECZnzGfXseU7lDlnHOg5JXbcw72cnjOeFBVNU
ZwZtr1KNv+rZtspJV7fnnfTyqc3dEIPzRAfh1eJtdSOG7e9cVmyN8sme/pG7la8KVLoejGRODZME
IgFq5HTbBu4210uf8rw48Zp4I5d81QbNgjkvVrbIiASg9IIcTSl3QP/7+KJ8BBFmJ6C2JfSs1PcI
eqz4G7+CyBahTa+V17wH+y/wjMIjXtVPTzyw6Pt4EU3RJIrcRh8vn6/rAUkoFI/4J82ZZO8ayeQy
Hy5mAd7uL6qVphFeRQCeJyM3quiH0Mksvojr3dELD0PJCzZym1ciGlJM1CwYhPlHnUYV1GuyR/jG
qqU36xdKmM72WAyVvFLXNdpsmiXxK3kO2fOykbcBdGVrlERq8RDzFxEc2yZiw9YIbtLs72RvUzU1
Jgm+EymcK22Jz0DsFF7K6yqHd1FAbqFkoEzZU7+49BsbbEaLK82ChTqhSRlXFWg6UNZOygNq52RI
IGOp04ZTY52TyUeVgrjs5l6z0aCxnXoeRVN0sJ4nbvWAgjLBkuJsQaNmbYrCKvWHmwJz0IX78eUn
dlq9LArbSvADBlLpVJrbypiyr+IBd3Qp/2xHrjlYOA2bxTW6ZwdGplRhKuaqpzWfTzcTOvPbp+g3
CmkuHerVio2hlti7R/6ckBhoYAbhQXxTxcwRyg6XQi+1hAqfQkzpY8oyzEAYcFu5kb75m8pDZ67L
Yu1X8IBwJQDPo0HFUHcScenwBrEatHbbmCX7jmL9lgQrxBF89sM9A4lnCC3DUNCPg1OLfR/rxcPq
grYO6KX6WDxCsa2zT+moNjB/lDd3jmRqs5SY/BpzkGSrjD2w/e2kDo+TkLU1bugStnGvWw1uRX9t
L0klddbG17RE+wLun5JZhMhQCBKgEEOIDMMZ70V4m7lGF1Hdlas4LHVrKn6NZyr+qKvtg4tm2wTU
oF5HXZ/bxQOt9Rb+Cunnj9nJdLXgtae1Xo7A2j1TNnfpadTgB0if5deA/fEz6BRf0UII5zDCNugo
qVERAecpUYpepvEGYR7s1s1RyObVz6klhIuguBhSY3jOEPRtfl0ePNrPrLec0x0Xa/LzFxBRgcSL
Mi7/gFdek7Lj27+pkn258yBs4q3ljQeOgg5xzGK0inufwPkxhAdnb5WgvAIpeI675/npIHct5hb9
OcKP4eCdAFDLnvxY9HCvPH1RI3PtuCOXM6sXg6bcIajKXXYqX2zWYxXJ1R0RFglQJi5Az5K5FqI8
P/EB/EJHnAXaGNVrloFiwLAIAvoX1hjssLeCCgJorjOZOLN+HlijbCaeTf0aqvDgC7hmFRyFtb0g
/+DmVNo/QP7IZGe8pqsVatFTVKStdGVYzJuel64OXZXjQK4NubrTrG0Yvd19XAr145nfV6X0NveA
E2Bheohk9LRmqQXWZbTq0NO+K1NAUP6zLZBL88m6qDkQQsqAVlTqsCLbj4SjbTZsBUoS1VBRpEse
waiWJOF0k9zERZOca2mzLEB5a/AtEDNjXlEVxskTW80Zi3YAMRY2vHg6znY/LBZeOs7Y1ZBwVxwI
cGxWlTYnaOe4Z9fjlPgNSQYrUdvqwMI71E3EsHJH1f3XoAqqY96nfjnh/QnxxjEsYEBRTVW9wAro
OKFV+9N0z7U84Fj8cnWo1rOqX+cIHv5VJERd2A0isJK4QSvmxefrYvXHmVXPLXGUxHsSvEqehfTn
uKARtDBNge2DtTc/1R3WOrFIhDq4Yi+4f2vi1x5l80hx5Xe8R+MnAKSn5lskGqqtlWLaY+AVy3Ro
CJ0PsppF++qk6asyhQ62Rs7pkKuD3uhs5WFqvSLaE95cqTXepIH0wrc6cggZgexr6CbgyFOkFF2B
QyOVIgCX+vkWafssfPeXlUShHtwDii4wgqk1+ZKX1/q+rsmu+kg+D8hbf5oK8wbxT3ekCDvuuUjq
g91JkTOv1ugKMZPnbRm8ijBqAT/nCwJUv9eUvgIIMe2HsgPAjz/jVro7f9Kpy6aiU+cp74aLRfc+
cRGWIVEhKBcUMLhAOLFtY28ZbCH1r3TE1eyYtAHfhj5CMlsFvYsGRnNpioD9IWLAAokbRGnIXToV
ClqDP/OYPe2GinzBypIPyxHAopo0acD/ybVCCXxWImHglWV4BQBnO+kPb4gieHRdpr578nl1hEG5
gkJ+EkMhaipDxQWBmiSa8TkE6sU1+UUUTurc3eD8BGDEtVsYZh9bFAVTms9XR822ZSmHFScW1HfB
MxS64WowDVkpcKTi7SCg/Pn+39LDjOegzxx/YRQnTR6vRrT2Tny69l6keRZLhOauhAIqZ0w6SP9d
W9yK6hcfwnEGNAlzy1u/OrZmTrn976Y91NtVCr3O8NrumPeEYrEffdMATJOdQWDneFzsYL49qmVk
JgfI/qq14YeDsL0/pR7fSOI/dhCAN1hnBFQibhGSf89en9RQGceL7ERRPZ9FCMv/EyHTFz5IEAty
Gko455w+PsWaum6petNFjRQrif4Stmalc6PZHfG9727E7SHrZjU876ddvF0cPbpZeyzEYHXe85Fu
N+GygohbMg8TsjFIDyGoM8PZUn1N41U0z7Tx9V3+iLZKWd6aqbOOH5bqduhqKgClkRP2V0Rs3/5t
ikb0NeQMfXdTm/uEKG3EtDkqQNQplHGe8Zd6WuG8M1k/Wtxf7Z5ac9ZC/2cTsS180I0J9EaGG+H1
u1oFtWYAg1fCu2eDtTOx/vUXWsEtgahubD5nxe3o0u1ReVEd1KOBL+XnnC1E8QExC/7jWfRKtyeC
0Erzc5g4Fn54bVgwaWatUgzCu7Ijb153D8XfrShJ/689bFClPcqsCurES+Sl6BOXMi8Qq9l67KV8
2lf8QsqEkFMRO5p1YmsXnI1stJeE2Pn3SEoP+uBXdRWubjsd6c7pp7m5oh/fO/JMMqHjOaXxITh8
/howBfdxPMr3g65YO6WCmpamzoh2kEU8H9OZixk335cZcisQXQ9Neko0HQFHJ1fdFVSE5GP1+O8M
BKzpdHSW/fSxpT4qmx/gq5uaJUtkw3MIHWpRzxPzLx//H0rl9lnAQZYwqWMDm7airoaX09yH9noS
+M2UnC1zcoUrQw6e502gM4v0nm9o7ib7yDoJ5g4zbI8TIfSVXdl4sKydFfs+1xQQsXq9ZenSr9sd
4nds9DbAp5ZtpFtsr1Ktpacjs23OInLZLIUolITZ/BP1Fd9JFtiz1j4rHYOO3+2+wsm6ts1nRQCT
YDySJNLlXEWXTVUlFYPPv9UirPqpcKPo5mOu2lSwxal9hkq41YDQLM0pWNG9YDuibINTxjpWzOip
z47DAxaAs75il0cpXhZqSD9KUDknbP02nXCBg28pOsOYLO7dRloUNFlqgyvMIxr1ibneMET3pvgn
ottxpwpeAYRSPx9VfXfr5Ky1eMSp3QP6WRqqK1GW0irmOGQzHVqzaRT7SwbkB5ZMA9Ni1SB3YonD
ZLkBZVxYHjetoUYabka+2U/6hK9t86+Pgy+fQd6caZnE/D0atHYkhBiGP1r2rOnM1VzCbEIsSID0
PHjpfPgedl2V2wMxq4FM01idz3nL2jn6ScJ/w1jJGmdjJuFOOicspdT60harBPmWDcLvvqClk813
ZAuacNlYaJfk10fy9BMLjTLEI4z9aE2GQ4GVQ1rST374vAvUT7+D6RLohjgHBXZsoPea0L3lKhDe
+o2K5HgBCCxoWs6hYK7tc4pAfFW3iUwrJOw3b4hjTPuc/nXoGZZL5oXCqp8vBXnq/myWda0I2TyS
BHsKrj+E4O4SM/mzQN7djt7i+rN5fCl02QKm6PhVHPP4OQ0ajvtWVthrmMjM27njLUWP4YSf4vxI
1jrrftGW2CC6GJasX5v6R8K4gz7Z4aMeVg+eLh7WG2NommMthJ3GN7FdwPtlYGeD+2AeuQv7Yfoi
a2NqaWanMLMwgyDX4TFK37WSEiArQA9oTJwiarRo5EGbGpeZwL+nl1crcLuI0Tbpvj1SaaNAJSyT
fg7S3pTUiKcEydvIv6IFlrWrtlTbQ7Ru317urburk8YJ/lIvsIIN7SprBSkUKENCSowcBijpiD9a
iDy9kymH9bWdw+JFn6y8MiMvqw6HePHFfG405pOibX7kl1JpIRydcz8z1Y/SFuhdJMzhsucijiLS
ShO0zOkj5GVAAx2U8vGSfrqSwVi7TM97LkA3JnWX4zYUMCb3BIEno2H+TTsEsXRxwqMyv5yqjrFk
7iCl8vb7Kscet9DUMScXgd9/YwJ2gRd3Jb7oF7n5jC8bZw7uv3XuXk0pAcgOgGl6omANCVjmGSWU
b81cxSHr3i+iIt7i5/ggL8M3ANygY7LqJOymEcydH1fOfdsevw3tOjmrEZKb+kwJGxfd2F9atrJ8
CrGWSv+EnfgPk0qVWJOLzSF+R2pWmUa7MpM1d/dDnqO0UUJbf3C/+J1jBaInV9dFq34qWagqhfpi
xBY5uFrmcd+h256GAjfZnozS5wDIZFLF7oE2/ACdfWnUGsctT53MvfamANVmE/OgAjD3OQxkEG3V
fIccYZkIS2Sk1CyYOXdf4/7IE66DOyPedSz07vcit69OJc0YUMCP9bB3pc4e5jakAIsPZb8l1vdd
dPWGJn37sHw4cKCKKwvbyspwDrAImCgLff3YFJ2AM3yPbmm5TY1+CGCUANGJ0pCPpW+RjhGRxkbO
l7DNfqtPbNWnt7IlJO2fsjLYYbt5gDOOEaW06qMbAqiB8Fbc9dTGRVy5J5QqpMxc9I+3geX72uPo
KF6Mr7TirHMF4l/4HQukS+yxk43xE33r/Xvm0Q0bhcjtranx8vjbZ+oMELAb3dVcAv9058Jdl1QR
OtRZV9HcMi0ABeOK/xvadrN734wrbtDYxY6Lf4vmRjIF/7Q9iuQKkv1upayR5b1NCBAL5a09svlF
sL3Roso4YDVx5bM+UUxBRBmlqzN9NFK4N0whBdcuQbgQhM+elAGgZYiPNKrq/dIslt6elCptMju0
k13ZwJmZrVDOGpmhGpJyNSPdBLba212fjixYxOWLssTMdaSO1K9NHXxoethSSX9fgpW3VQI8jC9f
nwuK4+DdHuSBQdlSTytpmLuhARqad+1WoIKsmvgkmyNPY2MER78BZeF7jK3rndRqazTpggrQGuPN
dx5eZIiZY2KtTsueYJEg4iBgSIaUD4SshVul6mbxUtU9Ei71PjDnPocPFoSCHScz9eeiCJwO9pjr
gSCl1zNtPKJed+iMfJGSpdorl721ZNYLYOBuDYMspfUwDaqTcwmUjBeasLxA0Tos127JM2uuz/Q6
/PC9sjtfmZK55h5IyjXsF347Zii8wBBL95ctUcC4lCRYtEnV8D7tt5gN2zywXYr8OvAjUEudXaeo
SLcujjfdGjKDWJ0pPZXMVrygRzvxX3aBa7/rPE+84ofuiGBsUD9z1z8Vi2oPCWanEXMlGcu0hpRs
0lrDg/unDL1VCrYT97SyZjG+aly8ipn1IAXCtYfZVogvYxO6XhzzEbwbIw0fUUdWEkmupLgQhS0n
ftrTSFY3KwXXNB5fEso8ijK82WPUwZhm4XggvYrz2O7N0yGC4tY7pPUfKFQnpVyS5n/iI3o+rhRd
0Z6TmtI4np2OaDu8dsBfxyPQo0eUxVHrVKa6dBzNSnMeQwyCPpY2LTarLqiceyhx5uelufUyR7ER
NVMjjYoDbHxWA/RHDKwCYNwFQ3RvHa2dypjtdEjVq7G591w8nWCdVIZVEeUbhi7z77vCKyt6QQAI
Jy1wMh67KxjlG7PGQuJpJ6DEULtRGNHCjRFq49b17lD2nKNLyY3jdYPM/LksyWAVaQ51bY/wh0p5
kT7zlDj4fwMeWTZeXtQcz13mJRCb8Y1UvF3FBbgkTYa72tb5XPwtEN9OCOwIPEm9ySs+QQfCDosP
w/uvgTAOb5EEhnq9f2mmGuLB9Y4W6cuwF9R5VmJn7ge5IAF2ftNPE60a4mgEXcVupTLLzZ+ZnxqX
X2QmpOSPELfGwxcAScdv6BGUax96p4en1hv2D1nez3CgNeUYxGH4yQ6X6Jt3mjHAQhuild2hgVyx
T/Mjrac/YAWwyY1APCy2iDx+MhP0FbxRfVN+r0sHiq3gZ1Xdwtkc+LYECUnEKLkd438Nmz0/DkSk
cRtrYJk3SMXLRdpkh0pKtVmK8UT1PUocr7V4amXyHjy+QLx9L8sGq4hXLX6ot8mLFYkuZKY6exwg
ygYFJfFGCLLX2oSl7nmqhHWCP7uGfZr2iwtd/d4JKWZusOIgUe9Ew1ytHMkYUh6bWXnLtCfbqdmf
ToDlHsAzchDmnblehuvTgP9R3BM6mQeWQTTMF7Uk/uZkdW1avT8BYncMJAn6tEO2rPKXSs6eUphu
nVw1xWipmwdNLOGCdil7I4uZMRJQSItpWFwTjrpqsKsPentmh0QCDce17+6paqBjsMORa27W33Iw
R8b7mWUvnxkqhlOpki2SrGW9Hiq2K937bOcqZYasQtAjab1i47QaPGeYTAKz6B37RIU9XlBVB8YI
K4RKpLxO8i2F8HjrGmy2cdkkxhVkVpg4SElqnBeMm1WVHIxvmmqU7VnSTNnmzeJsWQVpAwinga0S
P0cszLNYa/ED9Er9KuNrT9XjhJyRMC4n+x1/F17AgCcoScT3O3PqQe3dP9z3gLzPuzb0rWY+jxl8
4MlqmBapo0Ea64srm96+O6+gmSv8bhVaJC9qTBo6GLOtOhYUdHS2n3WxX+cdjGEMfDF4hBtYKRGv
mSfW3QUSifPcUbj5QXsTG58gaARJDDOI4Zgb9olcWEiR6S4lqZ4k1pV6GzwMryJv4Ti1bLKbpm9C
t2pvJokgMi6tgo/DXK51dVo5sBdJkKIT3OSb46CiDkQiUgnRa3Tqls30VO9BQwAeOV7Tkij8AtH0
IXpPmHAFDKSLkXuMx2lZHPgVzjkULEOYsbUKa2hXcc2dEWwAXBoU7ORt7kLO2nPW7nzgiaNwZRkP
JsIUCpNJJqNmHDrrHCG6RbcMlJZFKEdQFmRTrBgw30QkOMJtdm/9HwapYc+eTsfo+c7F+lFye5sC
mOsEWhqAZE+g+lpBzxR/BDJymlcXQXmacBUw7u8s57QnNfusxiY0oM5hmJIvROmFKEqdFkCdGovx
cX4vM+Wzb7cG9Efh4MyHHMO7TvYxSgsML08iWyTTRL8iyqqlpRDJ+0KRly0Uz6NdNm0LO7NAJTe1
6ebM78KgArHNklq6iVFXNbz+Y6xRw2HyVV8R03hlLVOfVqOIomsCYxNleZgy5yF9F3FpLcqS8zoh
B0Wu5OjqWV6DHcxdnNNqQIiniBQbcuJVNuN7xzimi45uLqaBKLgBAN/0ePnmEJoCbqSCAU78fRhM
QnLbTb1rhejdlbDR803RkPoKeLm785tGAATbpeW89tDYAdC7fl87TpxRu1EUiFskiAIw9BbwVHly
XMuzHzPWZIrIkX6NBbxT+0Dk2+hjo06GM1AVtyRPSa9LbuuI6St7L45dFR7giag8kgZIUyU9hga7
D9pWZba82fsFH+VLgKk9Zn1PVJ5eIvhPKnbnrRpKP3SsTosqfUcuzpQrXi7lqL5wYD6vbBnvIMfB
knR+HPO+bxaRKoEnn4a8/nlOPXczi5CsYxNuqpZCWXCBEc7NxeiewsXuyC0g9ZPNVR5yjP9RxE7m
412OcNhM7HLft+Bw3Qok0A2zkc0H76peEdW5oJ5ha/bkdVOTjAY2nE7xqa5XG+gA591N7enObVYo
+wt6D8+hjkLUlTDO5R/3qKrzET3/jLh9HMU76QYzX88DN4bmHOaM77/meezpyNfoGcmbANN/VOAa
2v5OBW+w+EvgM4jLjEVGRgmDgVj+C5AieG14hddOlEP3je3Bka7ha4EsP6efP2sMgUKx+9EP8PQ2
kz6IltVn9Y1ih8xyAHHnSLzkke5mhc5vh874+kv0BjBGuQyS08V1VvJLwCl/cXyB87UekuzUF1w+
ccm4GsNJuJcCxuPV3cWhtbmWORz6O0Hw7NCc3NlaUy0Osd33hkb83SgKdHNR5/alM5TsQglkNQy8
MRoBLZYH3TqsCJ8KguuPbl7uXSvEeRFrNBY0WpJ+RO5FvMO3MM8Crxdi+Jx9aSGTNhUf6XRiOHCx
GOSgPeS1o0JopPXV5365TRzTH3NDJaKr7biYzqXlhzfeBeEXKgbRmtc54OH3ArvwXeco/c99f0GI
xOZvG8VaxnVyTsUhyEHW+6C+ejGrw2j6i5O9s3LTY4v8Si92TtnR89uEP8SyLARfUcwSHuGSif/P
HAbgawWqWjow66ld+4jmElQEDboLrYelijNZQWIhuKgRS9o1nOOlNCwV+7YWHX+2DOO2ta+034ge
qp51lgYtwGxix1z5F3oo66EkkTUdsOKHz6JLfQ6GUTu2putkiw3n3jNdUAyQRLnf27G+2/J4Jeir
xFUFlpkFQI7YYuUvP5iN+EzOghx+/+nze35knMdkV+w3j/j07goMmy3Ca4z4g5TuAFOMCjtcRDwX
4FsqpwMdjVESXYLrf4qQf4rt4Gjw49Tm5jpdtYRWMfTVCeoEJKVMVLNf8GTPDv4DDXqD5srG/8Rk
3aYfT9oOYnUBvxEtjIjWP2qijalI9UXTUtJmWV6VBr+cgtcLwYHC1z69WrrsO+OdR83QdUawOk5C
3b8UCokJWCDsFyVSCZIMMkrgsGCrRPGLxGhwDVAQc93YytHIr6DIxopwbZdI/+pnu39UMedVihYC
Qq3SwfXZDisnI7zaOTYMg5oqdBIrHHb5MxsHIp2Dwf2fmuXdKTZStq/lAfEVfLopS1+wUcNVIi6i
OeUVz5vmoJ7GRiJnrZLcEfnq3vVTlqHVvYu883vTkbEC8o7g4VCzvzBqYk7nzlZi1x23j/rM4DC8
eK7nAZBuaK+v0AHwTYwhA63VvrodQ6mK9qemyLTDLOektpXB9D+4kfp9pgMA8+zHKXqun8mEy94X
W150txDK/mzs673xqlgfC2I2B0180i4ys8DJcrk/g8uKXQwjUviM8eKaiJlGsdSkO2ElshdlLZ3K
hvN7Vb3vFkJHQbDTPn7YdEEsrmPZensVoFEQgdJgrk3EHG10+RJXsStNwbXxnrD66JstxbMuukcq
ebHjH4PtBWc6nyCx2CedQNIDZtFl1kN9y50wDl2AAZqm7QKMvo4lF9fwsWo+nvPUCCGW3OATrXm/
E8AU7gL5IOTJ93x9Abk6quYug3MAliQEhEFQb1T8TzLI8hvueELg8jqCAlcNhpxkXK0z8qSVfEVq
hRPBrZsa4NWvgsJZLI3fsr4F9aCeJM/zouxbrA7Mc9K/tg0w+V72e1vOV0EpLUwsc7kNk/WSezWT
2J92L37hsh49a1cDD98d0eZ/Y6LzJfjpgjkfWwFtH3O3JYsuDoEmXmrsYsUwiFrvRlnCFBadyx+E
yH/rWfFA6WxGPTFphRIW2EP7G4TwbrXWalBr8/4UFfa5HTlHoKN55Vul3XkkgACXBWRQByHQxh0r
qvmXFgFq2tkeUofo6vT/axoxSN9wBUUbgp9qgL7XSgFtFnD89hzeDPJ56bR2f4a3aUHxYshXE6qX
dm/sOjA5120b544qbUfB/zDKXFKAxN5JAx42WydpIowkQCfr7ynYGfqntNE9gWksi9M4p7jucpKJ
C1//tA/NdEbdd2efN0iOsSAPu3P3kI1RMhx6wfr/Y74JjfuMgItZf8/jsH4pSOirhKO6OvazUHmQ
2JD9JTJKRUesKBEEIkBD8HzLNhUgPbPsmIK/FW2QKxUoUMcpjpNNZFejQYCcJhOBuKfIRodP6vSA
vZPpSVxBLCbYbfx3CSvjD5WdCUGyXBR/LqvfAXUZxq2g/QPEdEJwqia3JASEcn1cCIHfzKU9gu9A
ARkCr9pZgh7R/B+Ars/9fUdqvZdcf3ViKn/0pfaATISE1UznMmPwMuMrI35bDWrcBs7P92kiCWij
Zsunbwq2LaieXx30glhLKM3UPeBF63sajyo9GnBKnSeowBS2YxB/wLfOC3ZiqD3oJEdWMBHqADK3
PJxdK2m0ZCbJ2OOcvYMM1JE/2JdwT3y5twrhZwZ7MCLbTbPxhDEyTAj6zsxICtmEccV3WPPlmPgO
CAmG7oWmQpGEz7i7pr92fOYvYFbdQ2cqDp+WpInFIAE09uKeIyRqa7N663yza3gZQe3vhtA8FdDd
e+H2wIDDQrQGm+ZfgMfQ+L7ZKMoMx5t1HMnO76AVLBq17oI3wnDL8rr3bRFL8aTGwfJ1+/zqAeHM
RqAMG9IKbm3/Kr0/ok7a6HVzhrXDUl+P7OAs15hZsgnhuBlGkXffvJyJDA4xlTfIIC6t4xOfa1Km
7eoUx52M47DoT1XGLLenXXYTBogeUAtL2zCd12c/3mokT68qzch4ZCkyWpZUxs3hqDNE/R2g2Ct4
2SbTZERl0vZQ6xeh0foqdM/s1fB/Qxvl6FLm+bwkDUfz1JA4NXUWvp/uFNCRjqXuCkHsgJpGPDKP
e9W/ZodCfneDDorwrA8j5AdtN5FGPGhwV7mQK8z+taYeI3OMuf5B+1p694vClD2uvwjtR0KdSn7/
v41+WJ2WMb8keuGeI+heXNJvxYUzrg6CA+NBeu+Na32cDIHO+svFClu2rlrJqn9TX46zM++J+4xc
zohkixd1lrgj9STnhPZBqydGVseDbj1viNAtAF+/TFRRaZdF/LhrADHENF1WwcpvRoJrEZzSsps5
ejNEy8BOsfGAO0SsM9EW4/yPrbbmQ54Lp4Bj99RAe3SmnEKBk45wELmg6Sm1ISsg/XvfNERsxR0u
Z8Jyljx5yRkUo7HomVY6d8dcXJKgrRDr93zcoODZ3p2zHEnrDfM91Ywg0bGaeSxGXVnp0JCRYW4A
UZw0oNsSmVdeaJz7XwUhnpmxuJHNpw4tnO5qPmBwF9f0GlP+6txkx78pMHgQnAXLf20+Kn1Sml+C
lmk8CJ8bFtnini6uxJf95NiquoGsK7vZliGzS05KRSlilfHdPBqOBv6U4PWP1l7QI04/VzfGWNTj
HEJJDm/PSBp81rratWveu7LAYjLFf2T1KrOKFDx/HcDVYu2BwWFHRWngfsEmrHw6xeQUgwbc1GBO
i4SOMf7DAsG85AoLf3VKdrrv7S3zUp8WihrAO8rBgEjkVA67mw8dGbCXJFgd9pOsOXpJWEh1dgwS
SawZO8rnKWRtNXKh+dbB/cGyOCafMlGGEhKVQHVqf0TWVNXElHemD9K4H2Wpk5mBi2rdqvbCkdm+
Po9LdcREV56XDTf/HZcR0CM2xluThFZkhr3NirgsyDHjDxsU30Vt0gUUOkTT6u86kDh4kJT/TU2H
yRYj1zA/Ir1nlTX7us4vdR1NRctrkWGJuyWvzMB4nhZxrNJwsDYnwnZmMvKERuIQn5EasGS3H7GO
Ybhf5byAhYbrosAUna8hmDYx2G1WZmaGVqnJX6rMIFfzSMlYDlGV6RqUn+szw9xB0x1V+9d7dk0y
apbFqT/PKhNih0xMVUbThaO6LPyMiatnU7i75oPMHjSTUYSRRhrQoYib7BaRwVoV+xu2HA4ufzg4
aD6M4kHDU3Z0JWioNEYCUDruPMVEmmjGGRP6rGKj3RYpug0vKnzXNvv4qBnQtACfuek1r5GGN95P
lt2xBd74zI7HcMwr11kakcKVd85HszSm79yZ0iA05t0u9yRVz7s/TPbvuTb8HriBHXOhDLECarWD
chePtNz4Qh8jRcXs0gJnBFufjuYt9IZ9B2ZizNKq/N4KyGmol4bWaHqQjmrYizM2MeC3fuOCv9vo
4eER4ncuKq/FgSapKxfhDdojr8Y7thTa4Bm/AaWYwMBdVrhwC72AO2v07wIQqugj3ul2KSiZDbPp
A0JDKSBlBxmM/pVCBglLZL+D939m8rPdjMysACRyyfbb0gabvCSdiwcOljwCAVOGgnfpJk/tDJEu
wHJ2ODDJZaX6QkvnkjZsH7CutmqvNJ5vPl6/T9hW9BbAKJjxQIrrvNmsGjtHYFVv3nUa85eimcIT
FgPXZ8og5s8gV99p2nrox+c7RdcH5PIqrvmoMoFWBR2kaTvM8C6+c3ZW8GnQeq57f9cNxn8nbiGY
PbHgdwFxC5Z7RwQFzE4K0Pn2RilNK5+Sltx9xfWHxHjwc2i+kWFUmEpLPcg35MUtjDpVf7+wGEKE
ovZzrgSismNiaX2sBAlKAylmqR0ozE5spk8MfCknY2+XgMO5CUFllrMlphCcPOdr/CoWFBvIoK73
jmeueCaZqi7AljVgaM/8zw3EDCe50P/tc1MCNymR9jnLlFvw1G1I/hzD4abX5ZlFEN2RtnkMCE4Q
uEUTckKby9v0uZBL/Sy6B/HLKs64TFNFy0fadPzJXO6P2OhpOv2TkOrncoWweTgUXGqmltda81PK
GX9ghtX/xJyktkmj4UpOaDgkXzmJ1G91vrvW1zI1H9ksuHjGLj48ZKghOhQ9hnhOGwGiDITKNSnp
0smKrL9mr1WKfdO+9mjOtKRtZtfGjV7zM5OpXCc35b42jjPQLnI8hkndEdMGZUgwBALhnD2WSuAs
qcGu90znZVkaiYOUhYBhYPrqEcGLZOcYw+ug1q50lCTKrmmanLe5bzxndIi+ELnk1BOHth3uHgh+
TgPsgf/Yx3rEjumV9eRk975vnGoMtzrnanY+3sQS5yzCOA1VWE4zoKi4egH4YITnor9PHeN0gCcg
T+z8oq2ROVukA4xFnkEamxrNySlEEk867Nw3vLt64c6Y8uNy+1qYV2NKdHRXOecvpqmB4rxZXIqf
sn5B/tqiNCBATFmrU7sUkFKmEOLvTr+ctq+54mwYN8HgnRyf6V7ufNPIA44XO8T6JnHD0SKSsXOc
kJekz9R2VpHmBNLxCF54Gvxi2o/qOwQ6GPT/Wk3LIQCIovcrwkCV/Khm4pPLWTpOnOvfkaZGalgo
h4alCDPyB+wHSdJZFWkAxb5ACh4RHCp+mFcG8kaGoB5R9Bdzx++R3LXf4xPbzm2mAKrN1pezo4ry
0pGyvO9CtPH1DOMFqnxWEEGJNt22uVYxtfUxG/oRGizzrmURXmGZhUOEJOJxFfi/XqvgBQluXbkx
y4/EjmlUlz3SqaOjEhsENjQQEc76joPMBW6dd2DNka70ryWv0B6xRFiPQcA7V7smtklTHjwGG/qT
focbnUBNFZuEe5Ov8BXhDX2qtpEAVyzM/yYVjbfqTx+orxj0w0DNhiVMXJ9I4quetEkKCCNR4dEu
nD8PSJdwcXVCZBOMUDOzHuZaNGbTfOlFzaP86238lOU1xa88IIZInlnw/vezdFBrcaK8dFXLb3mX
Gk9nus/At6QxFXEzHIrzGbAg1y2aiMDO4II9T86ldSp3UKA85VuoXNF1hPAuqMezcseaB04x7kHq
ZYVpE8p8Y+Huh61a9cxL7WOy3TcQ9wYEHiA4CUda0mQMCjfwqaTZ2uKWc6d0El/4n4TNtlnBDPsd
1b5gw/2oO9QQ+KWeAxPMKY0mMOe2P44Z4LKF3XnZQiqj0AFWst2IEz7zVL+YxH4ybIXKt6+uO5Zh
rrwUg4AOsxaqC4sOJVI7UzpPPGDG48jGKiwJ54NKWS/S6zEVByCTSg1UqnJBZJgY64i1E/ZDCPBJ
FY+Umk/7P7TRiFqy9PJScuXMVUBubvQmFjZcXwkB9BzZpXmYc91C/3kiC8P3qbapNKP1L+9aRn8q
/xF5rV2odGZBRzunPLKvB5zBXH2qgym1keu/25eulO0UYHXCcL3qZXEflxWCGufhIRkRgNiME4wi
mVChFuazG31zs261JojwoI5nX3COgb6GqxhrC+IPpWK7NAmrtEHPZTIcZkQY7WJlGo2oKC/SgHxo
LhOSQOKgeqmV/ib/ugBkVdnT+hXifebw7O0qffmhxKyxbTdsF7CiqcIbFdBZPUoSOMNXXQhiCrMo
7srf34FAQux5QdWW6whP97U45ZkYXjC0zaF2GFRtHBOQVQECdMDILg7SuVDqRfhqrH9OOimmqAWY
+ZB8fwEv5C95uVg0plkLPnLnWpve1kUVYiu8eK3rDDrAD08r4pmEAjF/Z7r3Ckz/BFjXt1TogSpQ
dXX60felZgHhnnKh/G5tmtrxmK1ZP2ZQOpns+InvbpIh8xMI5TLCDgB2hNrAqVgJsPCgrmaWbwsC
qOI8ZJuNrvCxznUhYgAJE2BjY4l6kSreXainCgKS5rCsS8TiyPuyAwfbHeRnGnyzxYVRIgNAltfK
CzexuxR3G3r/j6wvWfjGQwTT+YR/8IGpVxssnR66h9gLs5/2z0hPgvan2lr/JxezpSUXUJ0Q3g90
SrpLMQHkbyGTv//Jud3IGiTt7i5JYxxzaqcxTnbYPZZWuPlw4VBQ0K8lUzt04ijswgbCwzCQKeUh
IFDq3O21nWuhfRWA/KLBLtvx2hXoKxkl7IasuYlF4SM/bruaA/chEM5m3uKM/DKSwPfUsJ11N25K
uGvo0afXHAubVEowrXSppcU3hI9bAc04UPXdpD/iteKBUDrcZyl7ysLZF84MfQ1KndkINh7NVTGC
IPgaTlL6zwf6M8rrM2Z3XtHNKdTW2/j2K35z2Jthb3Yl3P2be6GS0PPi2mvHwhlp5qiDDqSbHx0z
y4uJBea8/Dpo9xAcz5GsF9WoLAzVwduok8tpLHys/Pu/utRakYvC34cgV+GE/1CUpVDR94Q9nPg2
w32IxemH5ZaGTTSMK0I6NXiyay1IAcqU5bTlYD9txh/v+1lxwqvMI/m5HgE2GPZCGuGal+ID/KWH
VOKiXy1z6TTDG5/CsMH7So4A1qYw4clU1W3ULsANhfzOnHtTIznBFWq8/qgXot0wZQuq6yzwkmnZ
0Gjyj4VihzLqVk9tI7UpJ7AQI53vTZV13pM3kkxc4ydfa9P89l8l/lQdwsV9hRz+yOcy0v83WwlG
hjOAK6V8lQIa6ssYTdGz3dV0AC29WITWPR5FISlLLlCTsG7KC/bn0Rr0DwQkp6pIdMZppC6iCvi3
14B5WkoCLykAT85o5Tgt5oQzqdBnIgb23MSDygc6p5eZKPthLqeLeEKBDrCB43zoNezG4t326K5B
wFLCWP6X9NK9g8SX1LZt3X1E75KawAwPhWsWFvHjR+XKhhDvQAus0ZfX9T4gunMidhf4uaTzUs/1
shWXLvVgrbPAxjQSPwnw5oIHhF2sUfIhhBLvze17EoEjrEYZhgJi8ErgEwm0EqBJoR6tSMd23/Eo
KvW6Ml8d+oroCKarjRcLwdDZSXQ5PNstjvHNSRTXLShsLq8/MndDuaYfGwi6k+ku19Y/56fZhVGW
xah6zE7mhRi2+ZZnQO87CJygzCP9kt13xKVA60E6A2Ltd3iMaxGzJV8EYTP3Wirfcu/uG9U9fa/o
SBg8trSBS3vFxLDRN8S4/c1QCSMXRsnqefUkCHAYOsuGJjCbG9XWX1ISwZrqb5NMUHlEo0erFexb
4wY7UoosVbEUvCTyYl0DZjxjTPOxY/wvbZQACjWRCtDuXdnJCKEDOVf8SQj9K8Cjzf1KposnDgd3
x2plVNfKAn0O2d2RtRluZYuZmhL3PxXIlYME+QTiJ04dLDAd1fz8S8BItUtGfLNip2/S3dTel0mw
hVzxMwaDdB4af/jlQScQlug9s17GCnAzStGEz7W9f440RWog0BO0pUtQ35+ei+Jx28mB+N2nLqkw
4aFzj1PNzLyxnVWztOysg1j+mIPqypgBEQfOGIFCrOpwEMiK2CzaWEIOVu0DWyVNlmvTgJ+5m8Sr
hq3IU2ZOkmS27jbvdvz6W0Y99vCT1570/p0IKtZ/aTPNCfh1bp9FWx+kMHlvX+sh0i14gIt3m2rf
SBJq+YR/EcHGktb3Kt0C09H/W+LvU2tEgke17ZGstcKR6igdDKl5O3uDe6Fts+TYmIWjLJFjV/jF
BT1RXm8M9Ivt+Eswd+TIWAJNeQM6o066d/mbrwrl27CwVp3vXJSbFKJkzEXGlI2Hg2vHgyFAbSG+
611kLeKIARdk5ShEgZLR6jMk/F0y485ZrMGG3FFHElN1CXCE7RCNFdtUWcCTRWSZJDabNkTCq1rO
zufCsm8Wsbcsbiwx1fV/5a7UPdcc/oRMkq3yWax40DID2AFpQa2eoZqHCEWZfDwTRdd0uA+WqY1Z
h7sv0rgtQlsK3hEles7QdUNjUKLT/BZzLdxYJ9QNYD48LLKm2fErl8/jJbw9AbscDkVTN9sjnf18
wLHhlretF18ftR2cxy9OC+fgbInosyqg4bresR8BD7slEj7a6AjOJytL4rIYAwjXPHd+7Cgib2/I
a4qgBblzTUyngKDdDegspF8gPLNLB/YXwYMBu8sUPDUVfRpjkQ1IRx2hchX4fT8RZhZeDuGNyNWo
sebokO2H7AmteoWezlrZtRuu24JfPjmpqaOwplTJx0FGOy0GEgKIxQKGLuGYWXHJLIYkzRFDwZfa
hskr6dwo2TsjFc8QNtF9snnhg5kVcvVdiN18oEa5HB4cFjSAtp02HtSxS4aUy8Lw1G9v0yJEhbD4
z0ZR/G3VTV0q3WLQgYPyoyHnfFggFx0xylVUR6rJlTsu52DdBvgz2P6iSAhAi4hbtHOopLX6ueIw
8alEO9AY1gXEq4HOguDqqY2pJDl/eTsXcGhBhWWnInxsp2LaIir70lQzcUr+yxIDi+wAr9xvYuwI
17YkXNGkYUkAfdWMZ4t3RJj7gO7S5GNt3ObWCSf45Sm+xqbzVsF40x6aAXlxuzqtlyvnz/VnIYQb
qrE89OMN6rRhyTeMHDfdXk28q6EEKue3snmGERaGmCkcKfe/7XoR+cvjwtcrQJ4a5+5qT7H7oUmV
4UjVG/LG7obEVbNDwvW9/JhXzP3BNEZF7HlweHnP9rLit0VRq+8LG8zPiphylfnhl1CLtx4qBkCy
NI9gCSsZ/bTHfAGL4s8/E8HSA7oAjYT4WOK84sErw8ls86XL360OGHpmbQwykKbDFLepUCbrI0E0
ApBnvgCz2rbfBg2XFcobd6QaJ/VvPsCwUSRGt8yN6niaCnEny1CZhZrR0xq1ZKdyG7K4oEYk8WeJ
RobiCk9b2+MqTgTz8qwXPrQAkGWoiHeCxXeSauv3DF+YfpnRbmrg86Fs9eow+SCJOaAq8jMeGuQR
uEuYNIbEXd5SdQr5MKhtxwjDN2Yq++ITKwGTgI32ZEzlFeOS1UNkEInuJiEJR/B6NQjHpF1brX0A
U++EPSnx31A7sWruTGZqHWbr4Q9m8d5FE+6gRAFth3VpegaaN6EHD3qygejzzJxTN86MNNODFr7j
6jD5GxGQiVf9FE1wAyQVsdHNh5elW532X9kQTBe5uHVWLbEHmiXdq1dPlEWjXJI3Hytq05nYDUow
ri4QYv8v/OqkJ6AvOcQwh69tybIHxH/wGnz4Z2ffFBEDILobta2meTQBwXLMYk/nUXlwEodwzjb+
9/s2FWFwHSccAWxHtXd2tUMmc+rI1s9MEUiBHA+BKPV9L5D8te/xKMk7SjMIQ+Hq6XXiZJRU7Bqe
K1LWizZEWLtS4JEb1VNcshYjU0MXk6f0UEWxolkwoZdcVozvsePNsi3+pIsgjI28BJzr93ok389H
totpuq4DAyS7GES+Hp0WyNDEW6ekINP2vGScl0nkD53zKofuGhAeLR4XYeP0YCWmTmDhNjoTSe7h
t+qexR50pKNEnOwnXcYZof2uLYVxhK/c8FDh8dqxMd+daJOukTw2omNLMK43fcX5/N+wZBNbyLL7
YQmQb306M0xnlhSHvY+Ta6TfoyaSHPE2qzqeahJVTQSGSTHQu3DjSr384rEWjrpA+Bs+fgygiYPi
Ow2xuZsILhuabH8WWzwf/vqqOO4/o4jHkznrdvgjkaxdHWmkCWMPCIaFpzoo2yefXz1g6kz6GAA3
r2WrH6aZ1OyUYOiPF6mi3/9AguFncsLZx2MeCk35lQvqv2S5wlderKVC6lovTwxRfPJ74RHzciNM
1SJYwwyJ/EYUglX+S3Gy7pqnA8KmOI2Vq3jLlhZXaNxhyaWKBgHtuXaA85Uf/Y9Ee9zRISiN9OJ9
3ry8EPU7o/jjt5qUb4zaQIwvwqSsfqLpV1iJ62t2og4hMExFM68jS749RjT2jqCX0RyOgG2vcMP1
FVSBVSqd4ACXOpImUW3oymQfrYaMLL5DsZHUWbM1xJakcLwyGTTs7JSxcIu3tE/+9HX5JvyYuqv7
V56HLHFFG4IAVy198GMHEUgYz+hx3D/2uz/QWWk5SXnrc9i9mAPqzOD/vzWlGVzYqXapyBe/2yF2
25YW06XrzlkTqxOhfu8CD+muoEQIJ/BEAghT2B7bXtD7ewHjOywpl+x4eB8v2h+/ICYKRdoHTjAZ
QDKeIfwbmAXLStU7/N2v8aaUrQgeHaNjWdwr+9l/+55gm9LCGG9fBGCUCGZFiR/8G99hv1e3RvPE
VJdUDD4jf215ariswu+CCchEKoNmhZeNuvg31z0IVSjIenAr9a8ttZz22pivMTn5DGMPe/nLIbF1
v+MD013A2tPl7c2dnZW6zEBlkT4ZihRyY11Tn8RIdMGF6ncJQXFBUouwGUKNBwKKXrxLzpdGfJkZ
zhA/M8a7W6s5a5kGqxMbzd15kkXeS2Cvnhpw/pH52r+X6/QzmhTMmHUxDtts5h5uOd9uEKVRlL4c
H4OYVQ8pBAS2J8jP1Bxw/qt4zcW0DGJL0xSf7GQftKkCKTXSujPQZEXOZ0vsLHHo9mjc8zIrvVQ5
F7USXAIJ5s/ALMmtl7S9C2qvjHyaA5BCIY2F+RXLLsYAisN3rxk91OD5MevTjQw87BYzqbPO2p5i
QtzJ3zZlO3ZuNdPpg32ic+39vlt+UXE07k5vb66QFQZCd0hPsC/1oAx77yU/i7PPYsXrekk5wtWX
WqxrP0JWgph0x8qWdU0F7n2R/znSX4QNUJA0bSWcbOHUw16X68pKgqNmT5k5stDYgiLRrCR/wrUQ
wZBBLbmhRrvA6OXLQckYdjRvdEro0f7sFa7l6sX6Dt6tIKTvbcLCN22z9OVvWKUhOsyJFwfeaJGL
t9EMEBIKXVlemuznCkwM4/DQBa+b8AT1FWl5HQ1ffrb/M5OPiIdMj6o3dv4ZlCJAhMfsjnor1w2O
LK5jvMHoiAfeVDHH6VGVE4zyRDh65K4h3KVNHYj1/ZDyNYGiBWFQr3l7WpT0SxNK07Ldw0GofQqk
FHV1IjaUumI/8fBMw4NVnkAiQCs04jJI0aJwjad9v9yOB4lf3g7XMomtooKEIuOnVH7AI6X8tRsP
3KtWrvC8dqtrFYp+AoT3ZZ9+DXiFJ18atuZ93KOKDnLcAcFnV3ysA9W//wJur/u+lRrwep32l0eb
7oc2l4GHa2aze9sbSfUPATLc6vgitvYaSPjGokdbYfTgiULFz7NHxCLMAXvTQfDn0rfbHrzQsCgq
3lumtWb8Fme0BAFQJ7sC0N3CB9E3Pwgr+M+OBA6/9Q3wcL7oNCbiPoPGwYpqkfTqqoWF6mlzP0BZ
svUpTgtyoI+V17SbMfZi/qH4pwCYzNlyu+P0g49urCPOmZfEVSicPr/OJ6JNK+LbmRsmCVYv9zuk
38dXVcDhTIo09qjfk9B4dWxHDzxXim3C1fa8N/opAUZGVZEVpvjL7+aJRPvPs+ErwfNm59RvV3eT
dKrQD4s3f7VENnl7YdY7a5Ih7TxXnUFr9Tmy0ItoWtHcYLKBPJqEoU64l8LSpWG2NHaHI/46mCwo
oLXxTJ1Wz5BTXuo1Cgz13Fj2lyHw1wxfNfdL/qfZBnSe9uffYiMO4M4Q45YXibq1dUQfSW2UYu4s
7xe9Ji0d1s2fdV+Z4LNixF6gPZGLT2B58thEe5pviKnx8sBcxDjo1nF39mpW0v8rc+PgJ170s/hw
bsoG0sbGsfqSbdUCcOtAuv0ABpDlHLK3yQkVajc7gO75ACTZdlnVIQKP63oBdmFJYOfCwTzMpoYP
OCn/vSSl6I2BV9UlAWLEx4oq69DLXkqd71ZSNbSH3UwbF/GvemvJLNCc1V1GbWZgEVH0g5zdk3zy
825ap6+cAFy5vywAjhvLXFikWKGzkJTXyTAalnLR/lWBt63Gb+Kf5uehfy7Y+03l/UxvIXabb4S3
Vjx2Hrgdylx/5B4y22uu0FXBvFCBwFFWzrtmP98P1Ep2+jCuqivoAwo+mhHLeaKCq5p6RTy90Mqs
xZhBViOH0jC8cZq0Pr8lWZy0QSiJagt7umS48+prEkTQSoFPJCAkGpG55YurFu1Jjt32/toR/I0p
amgxmIrDH6WBhdxEun7v/foqLpHcd//Xf0BYDY0UCK1ThQhz4A1MnfeYT2PsmigrhmfbvPK/Akfi
tPS5d8H9LCxUkNGRae0v7J/61axU3zwBCTNpURtHloQv6cFgG0qnd7uF8WfhCNrVEe8J+4lxASPA
DyI1dNO5qAKAF9C5odMh4TLilKCj8cFThz6+q3Nh+24DFLFS58LOe4918YvNgh1g+vgD/QUCPe1d
PK4Piy8KozXMkD5hADCkk6UwDUFvsxbpnAcpWXoSZzZwqF7sIIMWxe73ZwIo1yXqVt2dMCn9mSeT
kS3/XS+4lxVWOMUaeb4RuPtJ7fQuZgKAXtDiMSkl6j9ZSAs0kK5cEo8tN9U6HW+WucJqyuTOD++Q
xG9bD3DRvh91evB4BUVYsnDWPC6gMkBpRI2livaH26ib+K372sOvBYRaCDXdMb6gxt/ojHLzneiu
mP+Yn9c18pICI7rgwGOs0N7Keu6EUP7gbwn5jDyewgPIS5rUUlofaosx3YhPmcyM1LFB6nTf4dQB
dhtfiiHOE+BddkLLcScBKZqjr63e2HTNrcVu74qjn0C9nSFKGc0KXr2W1qua2Wx76R3gOMpzNeyt
ZBxpRuOtitTv3Hf9keFhavJ/Y+RHXplGmPMoKNiZE+Ds6JcFiN7s8qRGfwbHT5kN7FMd0zLMC7cH
cWdFGjg9hGPbUvo5cCio476xrAchHjdLsLAcOOH3CKeg1GUcvozwpIn3UsvgoJag+QtrkvD/qjdu
p8QhkK0S2H8Y/E3/vOzJkP4swqA7JvJ8NDHCURetFyHm9vzaKfzpE8y78J2+tC3W1/bFwblGME91
XHWtGy6xwnvWmbHI3ahUOZd6YzzUYJLztydc3OqUvqD0lr4k8tXN2j9pjDCAeZzZT4ol8MeLJc2j
efxD+j0Ik2/mjZQdoVrSkTjJ2fwCbEo3NrUpxUYjYyo2pz7jtensG2NzZElyhluCVfWHizXgsu+s
E8c3SQrM4ZZIBJG46w9xt/q4ArpLSvX/7vwEoJWX7sQ4h29YG2Faav98xTxh1pugTqpxmyFcfwce
0NuVZ7420fXfSdpXs3bHKj3BkqmaJli95P2ZBZcScqDCllYXBs2f+2T9KaTsh6T1EimidT+PnNVp
Vf3S2JgE0Bhsry6jQUoU/i/rLkvE8Wsvn34FfSUtqvHieJ6dcf6jRjzJOZ7+fTU1+APQpXVq/yPW
EgnNWEnRWv4f9/QiuCSR7KKS+RrxQbjgBKLJ4gl/oRy165pO0i7nGItq/AVtqBYHUgzQPgQ43Lc9
RoOuaP3z/pm/q0Bi22NuTIO05iN5HpZsErvUAf/Wipq7X7ibVLULS0DQYGAVENCjvOI65dZDxAu1
CXoeCSQmZhDyntzaIa2/17lpN+tuoxE2etbmwYbc3DvDvuUaAnXDXHDmhewleTay+/6uRs8WyA89
RdA+LTE/mgXHaiDgKTosOEpak+uok+XBoCCdilIOPL3MeeDeg+ZPFYOHFWStSMbzd12lAIPyUbGm
HNjKz+R9oTYkSveIMfStKQp4vohJhL/yzJLMeZMEgWkL4Z6jJlnTzuPMhG/sKQxFz0YEEn46eKIW
NdpSDFgyasmyX3nsclzLwPJRaVaqDqusNnNDoHO5T0bn6I3nViMzC3Ehy37Vlz0tNLPfLOaH7jpw
1WOnhVUOG6DtHoo3v3EP9Nuli4n4OdlKrsy0v9+Q6HVtxmfjpOlBCj3pBfhckDiYUogZi+gFGwi7
o26ZHHlzMDp8yCDV7n70xUhorNK53BbOf7bGKGWhmkEVbr0gEvj1o51yu84bEmJg6IawbkkkI5pV
yT71JtakugE0pKPK5kVgITDUaUylDTejSXmi31hs7qz8VAqiMeF7ZRgItHqsUj9YM/EJjx2tc/Dj
NqCTI9nEvEHSI56qAsBKEv/ORuwAJGv6+taDYr93HYOXnAU1Wy0ytY+F2d9ZimHwtuG6nSu9VgbK
Nc8guqqx1P9Vq+T/xr2KPr3RrRjJLefFsjbSmK/9xIYK1OuXzSJ4sXR331ozhKrNOyojvIf/lcZR
JX4Hr6kwZIkoqwOr16SHcq3f0b/Rto9/fCYLD4fMwihCkn+MvYT/q0Df1eG7qA3FYAoiLNBCK/MJ
JDmaeEnMpRZ8Ft5yrWXxlNkYnFyHAma6O80SF1+0g5fnlL+hq0ldpQqh5hNiX74mg9+jeEZmXD6h
3OWI8V6JChmkDA5rygtxI3eO6MeASRBtMi7zkbbEWPpmpCelB4Ksy7M3QSc74BcgT5mmh6dNPR05
1g/70LTLez4kCmt24wfgYwdrpEPZ7O/BmKRN1x6F2nIUU2N0nz6XdEOSrErjiBRwKuyw4Om/q/pC
nV3Ma8rYPm0K0wPZV8ttyBEaO/fjag/BeNvKIs0qeKCtFIidbiiGB6x5qUZSpAr0D8+p2IgiMZlW
k/mnXd5dAKcdVOdFMnQ/b9MFv79i5bKJvHouu/QRC3PkzQ4bv4OdCi8OU1OYriDxzkTl79iZ1Ysv
5n517IIncbDjc4jMqaBO1eq776NaScGX24c6AodE4AuBD7z6jOIWDKKchozhSvKhajUcDi/ce/9/
UmckebYVcKcmgSJBCl61OUP1H0ojxvmo+s80kwN/iZA+nZfL37lBYBHJWYL89xeOSeh117P0J+T4
O/2T2D9PUYOeijKlfDM3Msw6zlbrx26oIm5esLODkYu5EDJxLS7AqyphNBMjqMiKI9bV5rNoMBNp
4Gj6bfXziWrz9YUfaNp3+YB0FIqe2SqaixlD3PvazXeMr55Lfb1PNMBp3qS7/WO2YGophVQXyNK1
nqiLrfltrtQt4o47s63tDQLCqedmy6aNipN9P1fc5w+1llYIWP4rOS+LLvldnzccLbOUNrS39Tj/
eEtYlHsB4vTKJNRHMp+fWp3EAZP974SrNd8NcxTL/yKR3UAB5+cUBApKA+a7x2estGsEIR+wxIei
Ju/rSh3hAow7HPjHlJIDPJwWOpIrYOZzYc13oBvn8Ijvlt16c2AnRd9lkjwbRcNln2/doi8y7unr
I4ceQKcMY1IHnL/0Pf+8yVc5eVSB/yGT+YRo8Ux7vSACrkB1pE/kFd8hBaLPWQJ2WkhbfmStDiYU
BbZQMhvYWmYG0ccVtiTrWnjLt/UJR75hiNM1GZhKhq+ID/XRRgbO3Sy9iY3WrZG12e4ML9grGehk
blh8AbdKD68gG6RGSuNK8W6uhEw7omMC7DFGiXF+AiWYtQxa4ntFP+nbcU8ygXbjyD7i9tLZFgit
RMAlS8mR0ivHy28wgJGXI4AKEc3VjhI9MVfBfqfB6s59pTdLxgPJJbkUBIYTI3nG/kSGKEM/HXRY
9zvM5yLd+oPBpPqIxYjjG+waOCOzUwIv1ZgVizxgcJUTfNmoCE3F6nDkFR1C/RDMi5G0+BafIUGK
zxhZeutXhMUPOZ7CpYmYOkCB7O7J91pDWFEn9Bre5dxv6u9qaTAmS90SP/3TKSJmUkam8I8eDVTO
JP9KTdkfVSQzIJeKFz/VwcMCUQ2vNkdEXKqdX4d5XtNTfHdAn1U5UYMzkrGPJiCHhLd62QVeiMIF
iX84SEk2Zra1tL4NJ8J5zSWdjA6yghDUhLUYomSnIDSRLUu+DupoIIZxTj5qGNgvrNVsschH1shZ
3FIZfjgpXkXlvA+fmzeq9xwb5v3NQj93liyjWwHWcATkkuGFRFoTbG2b8dK6NnJCAyvvig5kQzMX
LPBFA5hCZvzIwcOSK+vqvxtMhCBpvfhbceu4GB8KF5z8zY8LCUUZWnIPzD3qUarfw6ZiTzedcU8S
N830bENYZ1DhMSJiDZ6Ul9QYTPLNiqnWZ0VG0da7H4oHBFqbc4Bu6CXko8zUWKtSEaar7ozxVuxn
F6izzkRojn5fOnClyDrlWHqizdPulA4DBOLyfXkOATJzDlu2lHaOVLwutgn/EoQk2FC+fCGxXkB8
XyYgGgRq8RO946SU77alVum+G2dwYyBdiIm4e/TAVOnLrVuST5XTTZKcMxTOrrS/GQ5cWDkQxmU5
NviFwuHmAHh+fyw+ucifKOAThR9xtEQd2dx9BlcGIte25k29CBD18A40VqjSl2yeO8Ihh57QHz5E
aClvW8R6P5z6+4D3Q5orv1qRjWekMxtRk4eT2ppD/C+SiuOnA7vRmr3uFYngn4yG0cTlSExMcH9O
sASpjo0g1vKvd/maY8NnkczNgZ+Np9XVIbYFA7k90+oOg6duVngJCjJ034o/JDIj6l7GjASxwApM
qj/DxWRPjBBL/aVUVJoNZz2qi6+QoMZoWojM+l2ZDaZRrRwrOgNgAP71tt+7BaWmSWY7nn8YsO+r
ViHJzFdlRWVpd+a6OwTHAgdulVSABx3g19l8jUn83vv5QGg5wyfy69YDxL2mncL5+fPT2f2JaTWS
GS5sSpr7vKTVaP0rZyPQnZghev6pmwHcCtaqhWMaldgZY/FiPtENymi4GFLj1OSV41LpKEuU+k28
5YH7ZvhMB7gWpcuzl6MNh27Vkhz3s+ziKVjXOkZ1Uebpk8ekrMYTaDYF10z5oXVMksZ6htsQ1QKO
bxv5AO6ANDfod01AoJ/Vv9kSEUforu+BakUeE2Q4ehMIopz5s50Dpg2G3DswvXW4b/AONZONPUNC
gGdX18oVPpZFyQeNXGqJvPyrGiWHO2lztgs1uggVCz0WGNuGzwP1N/ejLAVWygRpgI9HsFgtb33U
NpXdsrc2g8uebosMMkE6gzm5AiLUQJH/IvMqXGflLPhq/bD9MCwJdb+1T9pWaZ/xvwEPM1EJs5rB
EgFCHPjy28qfAATHTd497fk0HRg4leI5o28UpY/lrcd0cQ5Nu5fAFqBC7sKDbQXrhBc41QsLpqEt
WIEvPR1/EJDKbJMcC+9LWnT222Vd2JBzLhuxSUKLMwtrI2t++UNPRiK3xEcEE+uWjgO2yViMs2E4
rcAJaPluWNy5UwJrIRcPWEsIu6zJz7pms7+Fg58XOdsXtIXDIcoSDSB1lHmhxYc7S+9tx7pMSC3a
Oyvg5bzuGujhPEU9UcnSczYbeSzE+eyNPimCZWm9cJdCV9KNuILN31O/2iFf67lWWG4v1+iFvxmM
D2k4E/kJrQVC0lu+RweiCX5zoNItJFmIAJesi4kv37pRu8mvZm3Uviwu5SLhUv5ROrjvcW8mki3a
WP4rwifPvTiyrUlqe0JfLAiVWjx44HnmWtF5tM9Zd7JZyofnO8TmJFNuZIm7FjNMBvfYmfxO1NmW
9s8jYJgMdmu8C9yTakZ3A6xIVRGNbHTeUuBpewEv5T8VeJhT7QEP5hc/ASPo0P9+Y7NcOJWJPLBl
e69gq1G4saOEmRxU03wcAMm+t0Y/LVNNieSuHDjMmZpjeZr+f8tQiXKqQsoRVx2vePnh5SBHiiCa
YD63dpAhcB1YR+HwcrHF876MbKUsa8V10AowsLkVYaEDR0txb90GaEBKKNn6uqML26/Oen8Vnc6E
BpT21uUM9gUGxHrUcRzOI8qE3i6EkMlQkP2KWsbjD7dHaFH/cvp4fl7Tev9UeXp5pCtyg7MluEqP
u2ptHaJPShr1reJLtGhpx8ozCBW3k9Yhp8X9RO9em8lBT+ZrurUlBEKnb4QGZv542n770mC+QzKx
hGyaDfBnk3ndyjp0yLgoPxkpNCsb6sbnGF/+SGVCqYQNJteQjtblb6SeGfnlfwo240vKQXiHDvVy
po+pKmygG6B6oxjvE1OrGAVkbX8M/oBUd7vNw2PWbNOaQr5lFGQzyt48DZnZdMIfHtQeLc89G9Mh
Jg4vH1xTXOfEKUKA2E2jbChqPps12hi4LqzDmNgRDppwWvsVLgP9B1l1LJoFi51U611bSZrjXuPm
b5OXpjP6CXr/8KatQU+7/bZTlm5/9yqxXRSBvtx6t8wH/Q3NzbaGBLbEMFmCCuGyjy9yb1qH8idO
DKilYaZ9IeZM7IByh9xQG4SjjCsxM67m//LJEPkKg0MGzXambAN05xStPzugQ7ywlLLzD2n28e4t
qqb6irlClm3SdIfwwQ78adquAetCdaXm0C6NK/76pMsh/Ps+YkNGJHn8csezXTv+5pKVMDBu3wP7
vX0yEjZOCLzoT9valEVn95ulLBQKFUnaEBOIaIEN0yqnHL/sMpyEf83vzROYwuvtsq2CfUli3SLU
jAk060szkYiOLfGqCr90TtIN1u+kyqcR018Hkv8StLaPrqq6Ss1uXdCVssrP9ZKeb0laqu8HEigM
qwz2Zg51dkG5qXMSL0Ve8CP3RJNy/lARq5wbAEhnUuej1DfqkBAxQbO5UQ46SwZI7aTdk5bppnPG
2ycisls3fh29BkIonMGkPkPvIr/T/ip+2HPw3TeqxPwiyl0zNsDzr8tqiHNp+pQZZ9HGMkv/oAVM
6t+R5Ee0k37sP7UHjxhy1YGIMKNE4DdOc4Ch5ixiJPGrhfysvf7ZGa1TUj9nM3OC2P4bGGTzlPTs
vt43IU4mw04MEYgHmKnO3/oY0nFq5ruPnKwchkz1+C6U9UNj51F9b9M+BgqEA6zBjqc1cS5AmChC
KkQRZrIsg1br7eWBuir4hGESdflTKuq4G8Vvb+frOKZoQDhXWdYwth50YKfBjKsDJY+B70E69YpM
eMMgtxxlfIyuh3Z1vNJBtHsei10+oNUlrohEF1wOn+5KSoA9apgPMEYciBW8KUsEArvs3qcaUsLw
gGbAxJTdeuJFZ6iPKOD/RH7lnYuN2iCvBhPME55JwzRapDA2y/IJpby7o0jv1FNskNY+gofOuoTf
3bXeLU0awismf2uqSo5ysaYB3ZVJ/ESc98vcVJUWKfEV4SDhRKXHb6AQFeUBwbu4SizJMaHNCsOR
gFztvwNSghwbnivjedpYd2gX/h0cruiE74M4lz2o4XHz+cVGcoTGNiY06zYWJTAgx7P+s2S5e2jF
pTOCmZ8QeCpzqQvgEt+8tYyckjgSJ+ABDTzjRaCG7LU2oJTqCscB04+QbnAajQQiJS4TcMtynSeS
Yhq7lP7LFL5FVY/zlQwp608js3FVVNcU4ye0BiXGBzyIVTA+f0mgNpQ2m6AxUYGlXlFOtzM15MiD
+vnQjqhSzrCFnE1I70CXjCQ03r6Iow7MYP+WBCD1xZ5tvOMlCKH93c1cHWinWcEJ+lR4G7e8ey9b
stwjkdEAyLnCq/ei2WM4gKYKrGPNdxjGef5VrxsvnvUSPR9062Su+FivmQGIHbZc0IGeGWgXo3eH
wEG8PD+rkiMwKT9beJAby0qXs7pS0k9aX7x4VzoOkRu+vBX/xFMGLCONB0P2Au7eu2YKOwfIh5F+
2FAVRYVxZCW3hRntCPZd1HDqmTQGC6wMxplqtstc1BxvyaHjR/Yb9JU//LoaV/6P8UZHXhcc9gC8
XIvF4+mzO0SLw+gq29qrq+yjXsW1ByU5R/YUC8dDYQ5yfr1+xF6u+6f4UyYYpSneNZldEBaESMHO
OZc/aNQjbua4/u6z39naKXFLlAsxP37CWFSQDJu7pd+8UdcDKqkgcPDpeiH24W31pbiUKC6Vn0KR
Dog1zEa7yK7iOthcWDYHp41EDKBQFDOYicMaYcvQcaeRXA94LcJjTTJS7m9Bx52BNflhgWQSkmW2
H0vkEoSUDWmv5ILzVNtDM0OpHsRRHfIouVcdbCSqyr2xA+peHT8B8PJ6wpgJiInAW9KZGZ1wTYX0
JT2RvZBB5dVOvRYL/WQ/yUsgVkNvSR1Z6xdNZYh28i+s5BncIsU/XkyeryXASs0XazCStsiQ9X82
Vr8gmB3AgF4dZJaB2yA21cRtyYpQebZ/v4jA6AxNTDVOPtz/8U2Y9Ki4CB3N/Y+uPftcAcVXDh7e
2N9ZUWV8RAvZio6I2gUjcDWiU4LJ0fXqDfjAeZoZQsYNDLdhAVLdLuiMRlrsLl3fzq1nRcw7Q0p4
OMyRrJlUbGNhWTu7HvulAPUGR9uDck13fImWfnpmos+8wHYdpLqxAFA7JpjHUdoc24cEQvX3zXSh
Fubc7K4GlSMxOy0YIYDKTe8bTo11Ficy426I6cWYlY2mNO8D+oMkAiUj4ubW4qB9dEbnZkv0GnI2
IehL/f1afTaFLLUsoUhWcoARCvuVdmdV8RQwTjbkWlvaFwbXeNFTmaDkqvfH3uj8AVAiC5VCB0E4
9VRg/16cYHleM+OJxRRBwZf+rioYxVku4FJXpEn5m7HbJVL+oUXdrU4tCDfHh8bcoyPtPOnxiu9o
JvSt1bFXs/RBCDZyU2IMy9SnnVMhHZ8MAbMDg+0FTJQPB5t0NvscaUvi8xDPNEanB5fx4NM2SI7g
JNSwblz0JVplpzlfEzqWZNsVyR8P/gZmHYBmqXtUJr03BxkjD1R6JKyMowN72MdcIjf4g+HHQE/X
lc6JS986QWPl3+XjFZ5m/Cpzcwe/CieUtigh+znrRuZXJU5ecFPiUxWeU7CHnEzgvjYED+zIpJq/
YvLGD2Fa2mLotBgjm8F63ULSBhcTtN5wp2gcsHJhxEro+Fg6vDq2xQBxDHdn7g6jvTTfSN/Ghoaf
bpsWM9wanAOv9u8Ihr3fHPumtxHe/mxh2QX/gspbwozgFvWoloehaG8rRG/kzZxq1NKIi4f2Xgqf
92viUvDUg8eCSaqeO/eOharsIVWXH2SV+shPxl3jMcfkNVHcWumf3UX4h4KdObcFu2hKMc6r/f5J
f0XZ2hdnyGMVHmYVhSbhSxp58OCpjBStnwmqlCz0aOml7+veyPPCo5rsJYsQyCmoMfC72vfXk4UZ
Qw4aNmwGVb2lcIc99qzQMgQAYycKSNXAHYEwMbgUmKRaXfuIiaaC3n4/5o4whbOgcYjuQWBfwHVD
L/LZNZtKIY0oA6T0i8aRl7NUEyDx8BdUdiwhboTiBCLYdHLd5B6NRpCs1pWlzqMM9I5qOYv7RLQz
h66YKdIXaw07MRbncz8zHJCJ5yWKmL8mJ1SQPJY94n01kN9jQO4cmsFclNFVHMpubmMhnhGzv1XJ
iu/NHCsbk5+zuX0l21C0eL8B/ZVvoUQHLORCC+Wpmp1R7dPCdEoD/BJBL5wbUcR0ZcVAhWOlAbf7
1Am5d+8roFCHYwJiZW8wVNJ/9ciyAOIoIJFVmIKERlyZSBvO0NkEgV7JVpXgncy0Wq7PPMCws7EN
qI5xlPnmtuQLGycSt+cpL1dIB0CTaHQ7kaKXznhnbqWLZckAxocBZghTNj1AeSakUNv/AWKbMcu9
WesY1s+birh3mpGG5hIpl9B2GyTbopN2j/YjSFd/bnifHDnrVYFHD3uxL+i7a7bNiz1p/Bzh9k4I
QOr7V8TFqwRRxgr/DOJt7LVp3HKf7hKxli5eV9ZImKVzcaQeCgQaatsb/HtsSkYFqOefnRdXxp6X
Ca3kRFv2uDAIcpO8dyWWz1VQ5ffK6ApdjtvaWZRJB5hN/z7tpT2f3yTgosO7JrGxOb76YaR739az
SchuBwpP0y6imBpyFg7b3K72HJU3v7pWhGysXFsHjc7YdMTaemu6Z/6YvxNPxxOtVMzYkoieIp4S
DQRcnE0k20ruEJdpg6ClHSTRgATfJJBBxpB+ffk86epE5ayFETY3DM6fDib6JDjKioT6Me7+D22V
VHAKGqceby1u89thxNDC7zyOJ4cQJ03RaK8m/+OwCXX8E9eRb0OrdtSpbrcHG4IZ6FFPtriOUyWH
pQISc/PIszk9AQBYTV63KFF3H8FynNHYI4SNoxrjw7vekCzGYz8MeavZR9rD63Nwf4T5Ozlkn1k3
sXhbI0pRdk1geBQmwYtMtO3brBBZxghPA3jMvh8e/0lof2Tg0dF6b6+vmLEEcUYZyn0leK2gGn3F
Mr7qQNyTelsbXADDfEoGxSRNxm1V+Ed1e+7812fPT3jkF8tKr36yyVn3uV+9phqDKa+1abjfUuam
MFiAwXBi6X71U3cuPqchawyZnfMalVYa4klCm3oleoZKWvm/9eKsVjFTJ/H08HFBhnywzeyyxW2K
QU/qHpIuI6fKs1CBe/k28wSAt3gR0Zef90++3zTNwYLAOWZyChtI2aPWst7fl+3aM2/Oo1g27kke
cqPw8PFfBkDTCWWQ+zXaKNT2qhbMthDUN5gkds9JIrfcd1bfmM+OKBoaMSma/viUxrO05YHkFvyb
zkI8QLg04ghJdy8s3yMTVZxWt/du1j45sVATUXZSsnVZwjUbpVOx24ejsZnsp53kDIf7XztiBZYe
fYBnrkAl8k6Y1zKV0SJE9upL3ovggkdQrAktoqV4LlFWukE25U5egQHz/JJd5xhs9gy4Ef3wnTdC
bfojcjk+z3mRi2EVwjYu60D3u004kSQJ4qNPLYSc+h+UvQ+SK/oEfNQlEU/r+HjciZt+uDeb9fIa
je0dvKvlP5k/SxwwroEPD/xRELyPEdqfjyr5kwTqU5SvoTvLWHe09NMCw9Nxylt9ipvNvkHOnmg9
VXtwpoDc6K82Lqc0cu0Y4MIAS9sIS/RhbReYe1KGmBjmig/9/FaJBy532yh8Eh4ySK10M9CXaZlF
iqLzD6Bt/i9/a8Rg1Rv6jmZnY+Q3f12BZNPrqPpVzjEa4pBXxYc20U9xKchXjq6NlgsyrwNqcKab
SELnTmSAArDq4yiPYq8vj9qkvbKdrThK3icG7pponZKdDi1Se3sveFRt4o/XeRvP5ShIUhiMG2li
kTbxW+re1ImRgAFPZ/6qwAE1sOOh5PcFjL3f24VWWFrhx/WYOtKvZda9BemPGIF5Yn8Elpv5+x6d
tNOhVIa6Yq4sIHyHJXYhVCAvvbLKbO4R8l/Y7sMOgoJiUFD2RYaPn70Eshv2ljfct/gSirelIsk2
U4+9EaWNySrfrLJeXjI99SAxwX4UyBGGQI6Y3JWS5aMvhk5dL5AaDacBsDPIL3r/+XF+CObc5RmH
hXQnUbhPbw1ZCycRkQS7+wjtonUBgWMPPjDJO1GGFqtBnoQwmUqSdeoutGFTtGNCkEYB0zETvX+T
l/abuP5T+30FERTubS0vHWAxjESNUDDaClJIT5yIzRbffiauXz6hlorP9lAJuh2M3lEtciaXDj/K
OZeNH0nXdlpN7ugW2FlO1JQ6wTzXVj0uD2/UgciP3Doc2CIVe4ZOdDDEyXuyZMHx8OoFsV/gN1t6
gEJAtUTAWqodhZl/EGsGfbZYGP+B6VPhO5xLg3TSVTrUY1rnrVYnboTxkz1Z04M8wwWkY2xlwDyS
sDGoXRbeZFDKXEXl+N6beJIlsha2aX9YlwE66HNwGZ71FnVo2J8u/b0w4PAeoLpH64R5OLgLrTGK
pudqSxv5Gy0lXDXdWItrNp//fWxdbUGcx3H1gkb3MsaR882zxhxuQMmP2K9zzse4nmsnu4SZ6JVI
HTuJytN+rrvhF89P1z+y2ty00qGtN5SFhmKlS+ETsoHeyVBuuwY8R16s51ctyDNyOhzRsl/CAV6s
8cE4ZPmEdCGl69n4sdUqzzy6QpncnZzXu3jPSTY90DeyGJykzasU1s6F0dRBx/Rtkgua3fhWUCEX
1QfjunRkf5uA4GOp8nOVpvY/FtbsZc+uWDrRo3O6xSDQd3lxzys1j8LhqB0OwZr7z51czwseqUda
vEyPyCYWudLVJcRLoVfS/k+7w/DRQrDo0bs6A3zFNDvlpbuGT8BIU29IO/qf0jCxJdXOWPW8Wc3o
id2pwyUKQopyas0H77JvlEzx0buLtDfQv4wkgOB38i5nBdjpSj8RYKTPm3LPCx+XmNGvo5+dZCM5
Jw9lc2zCqYe2r6xb0CN7Q7rB7UcnzL8=
`protect end_protected
