-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fOO9BT26MmVRDtNkS3A3yjQHYcP+bHXZ+pTOC3f8keMB3htaz7Gq6kmwrUwQQSULJaglF/EJa/sE
Ry3kSySMDfkhF/XzevDFeCYg2gdg8u8uj6Xnyx5R2sHLFUAjxay6MsrKqsy3E5J/SByvlISWOqN8
z78RAy5uyD1fbGYZnY1i2hylwDJsdKLLbtefKeAGX9CeRfjP6OosinCWNXhCYyZqvBx3+GZnM2hZ
RiAaB2Iz9ghhl6QiiWWjlR8XybK4U2DWnFTLMWZjqWtkLrS0vEF9ZJMsm13lcW4TQp4w+VDBiEVr
Av4OMXx+VxlEVj9P1y7xWFc6Y7c9gAM5hHEAYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
hzKGoQOLUc4JkUaBckcsDvRZxVANwCh0Ho6UbACEmRoOQmX9GZSd7Se3G8eWfD3LrnrL9WfQ3v8y
YeP6ZCds0ijBp/vQGW7u9j1N8MkAgx9uwDMKs547JfEHJdsD8Vc2dK+sB6uicfzP9pgxge6rVL4U
6A07tcF0Svu2qFKKB6fESJKGwUnBpy8fvIuNpRNJA+Vr8xIjbVWIe5K2UPdDTkAwFVMTVGso95EO
vTLAEm4IIbVCQ/xcYeJ1ycTYqA66mPaBPOQ98DTeuc12StxXU0b5ZsevRsEM1ZDNVlQGftYlkGHx
IWr8U1G+QnagjMJpwI2H4upzOoDLz3Y4ArXfMW4WyCj+HEEQFnMjqGyyuFwV+5rLwhNfo3D1blIh
wblyEaaE08hbUDcmDj5skd0OMncR9KO1xlcXHi6XpiXRz8+elh+2p/iQVlBLcdsAV9RUEwZP+7N5
hkjXermNxXth3c+vQsceFoNaSIm4/Ox5BI3TIlHSUtheNEgzpSp4XUQSfXmfVMf1C+Mf16357BwU
q8RUTBgGKNb5fvVINEodF6+0hszkw+zXyVUt8igOUVZFrHm+HbVbh70IHiP9ZZtRB08VXg5qjHP1
InrUMiDap94e47xXh5/2KuzT+RR8sv2LBTnv8riBN5/IP04S0+W4cV6hZ8hHNpOAfuTnFvPGciYD
/64ijtK+lfHlzpOV2C3u+KqVbIKXZuxLfYNZOGqtpmoHY7UHwuQkAlq02KKTNtP9a4MRqkMWv2Uz
LninrIxdGD4dbUXsE3dFaSNO1Kkc9TyaxoRIYnZqCW5c6L4YN23ei1a5pwm5J9un1llUKJ5tkCE2
tV72Ja9UaislquMNGhmct7+LzmYkr2JFgrfg92EX1/3F4knHo16q1bH/EGBGXuKaSTCz83AmQY8o
uZlN7hIYlCiUrq4i4EGI9jezYbPx+pieOcdVv7cVLhQRhFReWHSK6q0kb7L3Aelrd3gR71jwUUq5
aiJNE3iBxrRSJ2zxBFjthZJgcWFW+J/uq9M7elTzL9nfzFo39LplTHvNVQm6nT4gtrQpNEeJfBMB
wmfZ9bB2T895Yzo0sT6kVmecU8o2g5AZ6jsFCkfH1ERS5LH1uJ3WFGDShWb5NhqS2uBoL2XKOO+U
IoCszwJ4dI6XSx2UMIls0puJ8iojKpL/JSITHeL7cSXt+arUQ5fz9oVr6aC0dimZb8yXtf6NgdVO
q+0D+w1JJ46S8t6miZeHilmE2mjmJLgOneZyyyIWSkYOHs/I9AdxVm6EpiaZxw+26sRFXm/gyXPN
aNwyzn07Yx4mYwFulcLlWWfXRw5SMjIbI5vSJuKwU/NVkesvYjoRDxQBR6OIO/eRnS2C6J6eW9zE
fQZ1LwDI+3DJY6q6n9fW6KjJPRxusUigosAUf7az18/qERcsSBKO6+r23aRaSJ+Vnz8D/1DPB9Tk
bMWzCMboeXFsuTKCl348Eikq7Pq7FKx7tbOMBCRF/bbnapbRafCCMdPZTh9gYQLe/GZYsUryazNE
+DHaCPwHAH+lsMfGkjZU0qUcvw5csVB6HMqbqty6CCw8WFzwHxLbh0mgJy0DrD+2MCmHrP2f30MS
+6tIBu/o7cFRdo6Nd+0kxxdMAgFN1XAQgyfr0PaFKUO5pGjVyj5AkzokR167jeqUxcUQzvfvIC4P
cFg7D97BlUUAopk0cbBLDzKYgKdSAn/n/NqJrZXQ07VDtDfeB3qetn0ZYKa+az6My467cbqbilfx
8PCR38ugHyyRVi5jqxYGXTNXCt1FqRlHeidAnX9zsT5Cb0iHEGGB+yRwy1Q/oxolA0a14ihh+WoP
RkZzdlz8nB+D6G8yKz7KkEDvYZ9ijv2nyd7dif2QXoV3CN7hxjus1ZFtWc4TjGCn8nXn2W5OMmZV
8HfuEPDEX5jWyRF5f87Q7RhV7lbSpW5rNjTXWguwwszHB1BC4Sz4Ycr0VyyujuqC4PHaCw5Z5nbJ
1O0cNY5hvBIl3r9lO4WByl4xs6w6mfd1kXEb3QjMwNhy/8YWsvvkEVEkaNe6DIAWntH1pMZenonc
YtwD/odyPukjtQQNA0ZfE21/aV+fRzRIf5nUcRAq4NMSod0lCm1w7hvS068v4p+dmYF3NTTDYnPE
tZRMHnEsmsXwVKy0avTlCWMXZz4lKzrYN4ey2vLpWa/5h9R2sAx7CG7MEGW+VT0BJFD7Q5XHwyiy
wBtwHSc4iG89vf3fjAEXkvP/CgEnspE9+RKEUryL3H0Ti0g3VedQ6wqCYHJi1rxB1L8K8ma3KpoA
Y5clPrBt304kTJ2krct9ScG/ZRUrob9k3Lz79CqkcCP0cbMpGfF2+LZZCzhcQlMaqC/sU5JNbjRc
RNeTQbP9Wd0VxbzEeNAZJLXgG/G/vC/El7UL973zk8djNXgrmVBMsq68GEWFgI+q1bgNhDAB26EB
rl3/bFtvX+e7HgH4LmenkrtxQBd+ZBdmcTgMTv0iDFmIzuOhh7PVvNq1tPSjlSXEpwpraHM4ifji
YgT9PyB8g3g6nOpcN9N3fvbKINW6u0Mx2WppagW/0iA3oPhZq/H2V+bWiMGYmc3cLxshKPRvHeL8
h6ObEUPittzOJJYple9invKnzUM7750BLtjOp09Sw39Q0z3mneeVRVTopFqkgRzUP9M5380vAXtD
f8baGNsENlZxNYMhrv0Yo2RbZSMlhe/VHnNHj/YBitGXLbfYfUyvHmekYivz4IH4qw20HoeQSgCa
r/ZUn53iuuC7r8cR+IRMTy7NFxSMWu7vMvyaISV6o2wXrsTFN7uuM/QxA0Uh2ZohBJsLZUmHueju
1v6j2nt7yvCxrWrbEQt6qMqOgIdVauSXAYagbQwQlgVYRvcy6Nolg1av8QqiCzUBPkhnRtYjbcK9
nO9UEAXzJIxbkIsI+dFCVMVQXF3FnFbDMiqxy5tnO0yspoAFFDVEZ1Hnyt+fa1txNQ76GC3zWi0V
2UI37WA5OlYZGHTsldRZtKGInCXld4MLLPtvg5Di0Nwk7af4vrOPqEeyaNHzr1vOaXUxmAjhc/hr
mZEB9VAu/4hv3WFxTXYXxbkvfYBlfQ/rnqyFh8hWWnvmDkTQQxLPyKvBkRTftjrlpYGv8iKHOwDr
ObcKlwsmNm0a0aN6OGzyp6/xzcCoGYxsFWuoJT6upC2xLk8flMukdZQruAfFHvjvMEi55bIWIBkV
ll4lpk6c5AXi4EzxOGuM+0E5yY1TRMvn+oLW9ZAbcpvhZH4XVOOu3QZQcbJdeM4sQR0p2QFkmaRQ
xrr/VbID0CTvNEAYnspY6IJqF2X7nE54vm8i4AgqyiM/xTwGys8MFovRbjQ0cl6GXy/acpc9IOJg
K5DwxXb3R/IWMNAeTnwUX6f4JPkAmo2wU3wNmqBwaT3V6LEEPAR09lO9kPt2ur1Qp4eZFGaBv2JR
ZsanQdCX+a9GTwY3f8b7H7xHAGaJFG2LK2oNekCnXROOPEDHZpMnq70uOdSGeFy7oeEU/OiB6/Id
7Iv8rncFHW/3psCBNuqbwUvp1nKq8rsiZXuvHyZ3dW+Txy6GCrjvCS3QiAaq7qSD/Wy9UeEczpEM
7D70hTLdTpVoy6RMeYxv6GO+byAFjanpxWVycM3dZ6RLybjOeQGPNNIWvrjLRPIhUmrrDD1QIS2D
TbSV9BFEgiewQEIJveEWxU9lyKPae0IIhBhm/99dvTAE+pfC22tw8vMEhlqQbEg7OPf8iachVp8z
yJj/UNn+Pm/0LYwCJaoBRjWWhwpMcIk3RVzL16LIuX1CG+QTo2Cdjbs47fkWklNGZFzlxdESRbVN
zgHscFvgGDCS3Kx9lBquqkQCft8PbEjai82FZuNrcb7vdFg4HGQwmKazLpmciGl3WN+ZIScbkn4Z
nioQX7MRjDObDZkWL0UeqPsjuqWGANYIUKAri9kpYSyqwqC7Tjgt4YEPp4a24CZn4MS1AUFRz+aZ
Rr04JD5yR7e8vpP4BqQc+3CKOAroTwoRLQEHXv1P0iWi6b4zCVQPNjpIFCNgPp78H5PJYbNPHdNw
JvKGi7NgNehpAVT3pyF92MDDFf22+6nLLnMszNH3fRJ/F1jfsJFMnUc5cGqMnw7h2wi0e/F9X0Lh
V27vYNOUleIsaUiuYA2dyBDcfPulue59PB0KnI1XuCSmu/rG/E7hMGFLBehhH8y83j0BVLum7pyA
tZZTrpKZyanCAmuaeXK6nq7du8bqGxC2jLckQSCRtDRD4fXhVDC8+YRlBj51Z68V88d3Yvk48p3g
BJ651tb3oDXCByElqEUIq3Jehbys7Yawq5qXkiD+P6s0wXZMIl2k0DgY5QXU0dF20UtQ8cQ+Q6K4
rXN8smfdWanHglpxCGiLLYTjlkrkAe4dGYUfCuVyT1nYOtXjzV4PXXR42XIRhefUcy0Jr+dJJxrM
1XpW80eQMdrYEv3iK3yivTqsnICk+gAnxlmfo6KysgKnirzvYlQgRAdqGqHFe5H1VoUe1tfA0nwr
MpJ+dusK/LgeuW2bQZ7LOCmazMRnDpIe/4YTE+XkXISiMvhAPCAFKaBmSdp/UHakl5HYMG610OM2
EI3662/gluHZwoVxO2RzOoF48V5vVMWdyyAGVhZCVkWfud1PM4KruP8sdzRMHlgg6z8wUDjRd+FO
MpC6Eoi8uP0RvfMDi1K59slayoE/Aqv4F/Bl/SmxXzytdotrTvOntsECojTj37kJAMcVk+XhFb/m
W50DGOX2UkNy6u6dOryhslZ6PnntkL20/TbGib2Q3R+9RnTiX1A+iBBDZMdUfvqSybJ53xl7XNFC
g9KBIG3wxYfTb0Ddzz2InPd60ceVtgTRyiL/L5WxgoFxP6iTHStWETeUG39Ft9I+7HO4b17JrRVi
uBXAFnebyUclelxHe3ZxkYX0mGYQaRFo9swKbr5wP/oMaDFbn2EMi+SJ7KZFrSpBwvGXVsg2dCyk
FYyDCcs/uir3fxWZLZUIbZJL1RiayvJ67RJax9eVg6LkSmqAnn9eqX654HxbZexrZx/xEnv/t4kM
IDI7vUSdkY74Cxdwzv62abJXKUt/J8+ZFSQZDHd0L88uDYS/G51KyP2BuH7ttAdmjUEVzi33g/tB
t+M0+pINt7tqRcMRJZCicyEcyDUUEM8DdZwN0cW5SQs64R8VGBFTyzLN+M085sQnvuZ/wzudRiJG
unrATEyiT+12ktUuFYapli1j2NkB/mwMB+HQL4DkhAJP78gT6g99LbwIJGIR3tI4AH7wUImMxwED
4fDlyDBdGNblMVwrgtMKhh77MGMh8jqWrI3/+aijH/m27p6s1pogOXWgT2hD6JsWouqNWMbRTfRa
JnjnP9+WH+apHxrvYedCLee0aT+SBRrqUkYA71ewa7shsycXvJxZiFqhq429UFmivEUT+TcasCU0
CGPtsRD50gAh0aYMFkFPvYa7OePChHMGZTDB0iCKbtZdsmlfrHoTzBlI/zk/ayMlNFcrWeH2nq5I
FIHTPi3U+eMVZNcY9zIAnmoyLTR19rWotLiHwPvtCu4njYAeHMT+3UcogKI3JzD/XA3jf58+HBap
9s2HBaaoed6lQ9cXFmcq0Ont9ltaO7rheZovh+lZu51Rts3nLsJ+KIwnfHp/MSJAPLgiQMuTkSdN
Q01vwl3hCDFuYnVehhHq0HK5S3vT+JSLd5P6gGgoHJRFLrWQC19wh/PDqcReIUATOlS4bZEHTbf+
rHkrHZy20IBqZLDlkTqX3/f+A7orqGn6sA7OyTHpmR4ev0yYGegdm1QdZ0cP+gGGMYjCDQveTrgM
lGUCUsnWitlCOktAGilxEb+/woZ7njqxQ6Ba1LFA/ERDdbQ9suH72xb4o6+eRLCyCaft8TaEvb7S
oiKnVdDTXpQqlbQjvv/L9zd+Z1xzqStIB8Qer0d57JzMt/5fLHtVN4FTHycuNH5tsu3MmLamaz4A
HuYHVFbUn6FXR2CiCZVZM/x554DW70aY//GFSB6Vd9/u5TcONz/rCapEMd4pgelsV8aPElcDe2vK
lTBI348xaHm5s6LcWnioI7fGr+nQIdwnVYSBcmEKvJevva24HGGaFt9/jqS4/2rf5yupMMbNVRVP
A/cwPt1zvgVX//Hp00nxDfIQdFWIxzmZNHKAGtIPK4ontWmk6hxxzqfJiqIB/wj+u/2aMwUWYq9G
nfLuQspwe43xxsRIQoPq06ynOoW2cagX7lFL7qzqolhKUttFNRuME6McI0L7kG7YYy0wBUjvZ9np
P+PAsinOuucpI797bUOa4YKEfHxoPoDxc+jvfYyVAWdN2Iv+KIkF+8JX0XGIc/gkRRuEbf6VS2pa
RbG/+2HUtyXPO/MaecNULfM7+ePvBlvjFSpUUzllMiP7yJDWDAKDDnheCuM4D7kXm90O7XUak36A
E4L2SAVdiOqy7TEfQA08wL4CdQQSKtQ3wvxzZynVKWxve8q0QqZjeWqhVEvJkiY8yih9nmEjRYh7
9ottf2VCYTia913CtTiFtuBKOFd6qOvGYVooUszcsvFycKYvwFYAUGGZihNhB9iDs7I5ekFJoaNP
jSHsOEL5T3/Oq2RJim2HUFWOuqhMTjov4KMAYLwExP9d+IRDpZMjrOXqRK4QTe9wvEwXf3VjaRzY
XFWAXixw6HIEjUdD+NDpfsTpdH3/g7bVoyOH1O4evw3FW+EYh2WQOriqPwbHk7oEeY5QsJkN18dr
MfmfmA98OXUtBK1CRxzxr/BBXa3w3NcmTPN/0puL4dHaaJucxqqJ53QZ/u56Ui+I7LzkjQJ5W2ur
8AgJGg9bLu0sK01693DTILRZMWryVMsVODHWNedHWp+MZNDCj6rsmqLtWNE2SASJCWjpe72a3euH
EyfR2PwVc5IOJIdOXNWYRlBTXGytoZBa1JjmehrqqS/wDTEKBDV0X4Hg3vNxxVXfqo6r3IdRfkxF
apZLpPRdmo9LSFQh3FcHaM8601akg9U13kLBPB+g1S0ZAusUpCNvkFRzket3kZzP3aMk9SW4eWK4
hfeTjqC9OphCyesyqIA3YYrwoGcDuOI8Wuq8cU/If78YFmyfrsisOYtPILGhOUGQ6bdgf2qj+ITp
U8V+dXAT2J8tTW6EDfXhCqkny12CR3FtpIepuw+qBjhw38Ka0FCmUePTwmvYjBtnOeVz0xYLTSjg
s+ri9jd+GrSxGLEf+7g1BIn+dnyBdnSYV0udYabqIWc2lqCiB8sYsS/eBGFwhmXEe7AuwXEMiM4R
y0jbX5la0bDljX+MxkPD6JNflTDgUx3AJ209cdkbilPtBGbVu17ma2BKbrtAaU9uJ65f245hQQjp
2l3g8pO3WjLbt2oyeZZdZ77cNaTxwTXwoKS1qWTSjLNYi7iTcq3eI0nHNlKvarKmxLNBuX5DnznD
RGkH+iILM2f51dXLQxCtEcQj3gvfWCYAA8ign6A1snAhblN7NC0XUym+Mi7tCHsVN4PeNH6XzJEF
8Hiq0zDoIwtmdq9g0BChGZUlLMl3lg3/QXx3na12NaOVlz2Rp9ydYEtzCzqO1nSjXVtCBNpCdsLG
oSVPVMK/L3RvAQy+r65Fm5SdIn8EE9cRiEwCsAq+Nhi8rdCZ5HPVd0LD7ZEeDmtJdUrES8InwaRd
+nq+fphaoJx12WFPVW4E73xMfwYSIYkfH2Rfli+Dg9bL2LiurkrBasEr4zBwFtSZSJiswL0ACMUp
neHJVwhIRS5/Oc3QSAC+eJe2Y6yaifmCSQOtzsKWFUq0DtI4fIX74y6Pw7QX9l3/+nPQ/Z6XHZ+i
T4FP8zCRQ9ybHhKl3prkIRRJg1gHfvInVCSxJTsPucdH4xVIVLQisVCthQrePEnw4QB9/ERfabSE
4xSLBbfaHgHYE1P9zV4Vnu0NXfg32hw1tZf8lzvKrGiS17jU1y1h3flnQE/ehIvDX2SchWQZfDYz
8ImGD1gGD/e3zI00N008Z06W/MkqFksZKD4gQntAszZJ1dBwXMrvmZtRnbfUYXXBbae7nTMxY/UL
ifZCGMeTRTk1W6OWOs+lA8k+FFGd+csLvuHejbPAt/8c3pSSiWonOg13fS8vv1eFESJ+cYhonenu
udHw4lfDpCxNOCSX2RjL+lJ1VcuAdrdnBM74EDV/pRn7fdwNYaQVAoo/F6JNp9fcWE0DyBCL+Ve4
XSx8mmzVWnkm2vJKbnyLiTroSJiKLK8kzaj3mWs05jindXLejkf8Rk7TUOVVqhCTMHVCsqr1fxtt
DwR70I9OJlAILveTxr1yop3aeQ8v+/F+ojNaNi/P21J7gwvu5k9e2XvmyzjQ8h9Cd8VHCH8jcMIH
4CPpoUSXScTV1ikqztrfBCb1dK4H0sScrB5lPJJSAZDlbRvwJAdd1tjTXM7q0hDpDLecgr+f5jPK
6OHgMegEivsSnGc5YB/tqaek9Vp8SVo9f0UvQNYJwZbkYFpQi6Y/xqey+0S0+UoQfc44X+8ktjo3
mUx92gih8NPi/iL9Cogesq9AVq+1xb0R79Jqp+I0jkrRAPKY7QBPrGwlFFF067WsfOZeTvfG4p29
NuUk8rr4p/xDamgkpqLHraH5Y0K/fQYUO4kDjXberrSEGzRoJ0izLWw3nZ8x5JjfS122Jh6iTpVw
W+yX8gtrBN5XNrI6kTJj0D7fixYzsDgvONP16qvHhFk8fTpX2ibJZx9cFGIPxhPDPq6espmoKjfJ
FuKrKiMEJBVRJKU9ukxbrPLBBSiZsHHEGyzX4XCExFyv8ju57MF4RKKWLyrXSN08kx6qg2pTSBjR
ycQPhKNXtCZggSC56+IDtWZPU0lRpy+F+K58kGSLkQ1wk56P0z1QNoW2Fj4AIG8blWY1fSnq773F
m9RtyJrQJLpHIprmqwnzt9Su17ZikxwhLCadooYpN9EvxoUetEdqd3d00ZULLLyUIQoaBb8DlKJr
Hp3AyseSzXcq/7t3X/eQhjl3abfrqDyrzF9lHGrBlvntUq4qXmea06q/BtPxsEzV0uRsFLG7A+d+
QHtz7O6uQ6keaCnZ1cOTqWn0CuXf6OScsGelF+ayWs6fzDPBMlrMWuS47vwIsGwevu8ZVcyXclRG
6DQE+D5lhW15gbzYZC762wZandnQNW9BgFioz6woAJZ0Hq3RHPuOZblqBSKHLkP0V2uLigXGcj5h
KqQo6rgrHt7vmI62cxxAW+Q+LPY8a/AlsiqLgigz+RCjU/M4VcwCKIDgE/bAGQGhWhut9xRqLzbL
nlWnv8Lv+XTqvd7C5jWfQlfE5sgNfDqh3myiKBeje/NnRSNc6pDIayd97JOdQy0NV8rAmxh4ZUCd
mz+Ez2qAmpdTfX0daLY4XoQ9RLj1HBncA5LZjwukF6Gp4/PR7U0OqRW0YlnNyPwcKj2hlDHb2Tyi
fz8WtskBWVoDsnEntx4NF9YLO2bbQDwr643G7Izh9C7fAyp5AsaDQ29ZOgspJC8BbTHEZHzDjupI
XMmYpqbA87fqt1jY8JVPDNIIr3KOgFzvuyOG0dME/NKrV+rXD7Pw4rfz0BgK1zKSCiSODaR9tVJw
fEIUmHI9rt4tGZi+9s0dAkrOl21nT1SNrNTljIzdO1ch1ZIzD3qnz1ax3Y+BBs16QxoXKrpFtFnn
h5itSioHUHZK5t3iE2ZMDDeOnRphgwKYTtYw/Hg8Rb+XwPKwnda45dPPkhmNxFHze9WekjfjVrQh
a8JXukhwKYvJrn6hzKQlV/NalyQrkpigTaFq6tDCALxMUK5D2obV2XGBS4ayFGca437maS1QJnmY
CNuCBk142jHYip6GOjDHIvNKF4rvPWDfMVh0SchpGBP9ya2fXDZu4UBP3XbeuUcpu53lRzm8mmtv
oLOR8R4D7T/OQ1FU9r/vR12rzo4mof0CdVXjPl33nLw4zkuhboesDftuYF8BF2VX4Z569pN7Tvnt
I6nGORHT/YgJ99IAR6PI0ivUh67qPVx88MenXZ3Lf2q30vV0v87XD8/MHQCmZvAYWPmtgD/bjyCe
wOXq7/t+hs3uDO6dkC0csAxXX0YIIoKdbu+aSQZb+pGcOPthxvdjLOrn0N8aH8vo1lVIoYiIDJ02
Xia5Inn/iXuzVPPnJTspALH6W4/5g8pR2PUBLOLxgTgtZ2qvserkSnDsIpMxPQBGMDDLGi3DmNb8
RneaA+f6gOm0thynzBs/yaQRPNRcJ3OROSF2Y3E/uy5M7yvYnLQwAVpghJgke8yxRdjO0YBeAUbC
x46NG1AvsMPx1VL/6EVFAE+xqizNXdarOtSBjfxwyDMGIMKrvUmjBVxsDdoFPg9y0EV1EYh54AO2
VCm3VMIPRpTpxF8mbs/7NWO6Ig3xYdp/lz5FrAnv4/WNNdTO3z0WmIzKcJi+PmryUzEVk1rtGn5V
qiRVI5KnccechKl+zEoSQBgx8i/2S25rJ3s8KEy3s1gqQ2MsCcZjcGi5l+xXfTuziDMewluSqA9Y
t96wzhE/CuhcnAg0w4MVicSv7K8VdFL2GG69+NWHVIfZtSAeuvw5BfUorKSSvKlR9ZjgHwrs3X9K
xipxTosqBv6JZ2FOJw8GP4fo5hCOoyMcjNVB9Wo2FxkDXlUS46FIM2oxPqIZMaOnocSbAmHOV7Ix
GspJGxaeT3l/hgg9uhR+ChxjBoGk9ZsmSC51uGzKBx4MKE5VxO4yna81iZuaOjUlGE9cdKuxijeo
BQ4OOI5QeWU1l6nQ3jVHFsgrBUzJQP2Q24cpi2uuKSEj1HLzXcwyesfG4wmnPL0OuNfTvLwV9DDZ
8JgZffhHTtUu8WTcU1Stv7WqDEC+osdf5KRbS4cKzDTF8WXO3NVFTgTHZnSy7UQmMug4+1HJZVat
0NKEcz8ABU7zo3gxb0pMFLeQhVulxwS3tGEOa+TW80PB6hvelHXh9blVogw1R2ieRkQjXTD/E4uW
9ydP28vNNjsaFSiYtdasxE9zqwsYRZ2c/YadinTgK05ujsITfCPOAjnXUDJVFZmlKQPE/HpwqaAu
GsVvKgqQT/7JvIsNJzHmHXYf6hJyyK7shsBvsu3REIAFTWDsicXFEunDZaPXCYrfrUJrdVK43m3G
Tt3UHaQMeeEQ7vOi0okWqHHk8oqKOGjc/oC23pqWPd1FVgjoeytEb6KoDh1KRWAS2PhMnsAyvj3o
JG3t2bJTgZR1zaiR9Hr/mi5lVLH1Ds/jTC7hYe0MWgFFj0DMsac335xenn3B4uQtVFnxtbJ7Zv+p
t7JZlmvFgnM0XYuUoKfdi23OxrZIDA7gtALnqN4ncHbgptulVqbVw+uvh4ICheKKaJxwrZN6Vu9D
xN94MWJAuHIb3Kn5oRz3JM4qexwISu8T79Xezmbh+htRMZJHbcX4HQWkQSS0yU5fzL/oApelnwSg
b9ZwvuzJwLnrjF0EIGQPTjlFMS22MfuaTDxZ1ThwiDicUxe2mYVWQ65Oaz00aXbzS6NCZTBfHgZW
xza3oIiwYynQewEnSOlDpIR8lgUEAjo5Tq1tVit5ZpdyBv78dd3YQ7QchBKdNiPgmReU7kPxXWlx
mKxofBX+blRWXH8wyfqN1D5x2kNwrQRng+pP0TOBl/dZhgnbA+dbZuZr5xlnZGlP6B1kV5sL6PyZ
q4QaNiJBziQy9Wu+jAM/l7UnUR/54y2K2UxkIEDsdTOEw28OlyNE6IWPL7HBQWSxLhE3gAHYzmQv
voMd8ii1nfj/MRPWmphPDLQcr4GXNhasXsulmGXFsA2t/2cpD7UT/5PdfuSSYDP4nqCotU516hoT
0EzWi3l0a+mE7aGn+ErHoyYDw01pP7mluLTjErue1JS0oKTjUqiFFKv5BiKJkzFH6a65w2QsaOq+
uF1+IjW5ll2kcwzcnNFeYEkSG5wUqtxaOZ0WjOSCU1vZlKs2YacrGs+f/mEARcP/PLHk/KDyjfMr
45yQsfUKPc19VpHohpjfppb9qekfrrl4tjnmBKlTobRZTJ7vumW5D9lggQha8EKtlbQLF2vXRb+s
BZtYy2OuPlrAPgRC5lK71MV6dtYM4r2mFyjPig9e081z52btgRWGm0CZhwuBUD8kBx3d7Tfl3n7i
vim7tNNNPDk/WCkSPuk9+DQPD0rcpO1vQQ7HdDrb77cESW8UCu2MR/eLG/wshLOf0Ibyu+FYXzsC
1rutADqoqKi+JobDP/ACUd91d9fNbeCxQGsrKdMQV45BRf40xz47sLj/AvvI/QRw8TkImgD2pc+O
xrQXWXFCkNyTKqCy04GUk3u42fLiCTxCT1SUC1pOxtE6YG34t+7YmS6J1FVn+8XYCV8dmJOeZ/kW
a7hiufU8SUbbvcgQWuXy7pGr7f28DXHX8bOcGU7M57DGzu7MdOTlOtYMGA9aLsXZENncJOKsiVPD
ik4rD+weJs4Ov5F6csM7ea9fd1GvvY2INbh6z6wJBnK4AUwIrh8RjuK2ZuVrzNhflRm2yxAbLJNh
7i7x7gu+K2lvkKaWJL3eeAtI01E4Q/6eJtPCRCzzq8v6fNJ5vuqzGUweWbQIreU7bhoWee7DIRhf
j0wkGaEiAYRsWytJvKgs0tyLB6d37lofLHAsp9cHkf+I0eZVeISOWpWrYVYW/tntsqbDPAh4Rloh
SbtV0yboIi/zuTeGhIJKkhZv4jvr6Y54AX4Wj2jZWmcWATmV0W+5SOacvtFDs3sHp7iwGX3FN7sh
Oml5ZPo23DV5gtunCO0uI4Wlesifd8upvnEjqJphTffDieDlp7z/LaWX+bj82g6XKbacGjvQmdkL
tiIJdzkpmQgOk8XYNP4pocHP/5FHhJXdnn4xNNoS0gHQXcoF8BCIpCd99VHEe5ZBg3yvXKIHdQlG
hlGZECDh7XmBTEazOfD1r8oZXQaitqdZLDrssvWhhGYVTWPtkwg4BStxxXovp0EgRRSYVC4RGLRY
JqkZOHDdO9mJEvvx66GyOMs+teHzyUIVrC5gZdMTxhkQTq4J4/y3yOQlKAstGgHyrBebPy4Fh/gk
hPgxQdA4d+u47pPzV8zG0kiB4m0NdfJwmzO0+DI5ugO+pRQLyyP0DegjpXOW+Ju11WUDtDrjXsia
0tdhga+g+vZm5+Z2hnLdA/7NhDKMunPiUi6G2uZ/XJQmv1ATOTC6NrVwCwo9A7/hBuF1OjsANzyO
i2nxyCM/jMn+LKr3f6gTNVpEiOSo4Vf6nPMTgAnJj+NmL22xkgxH9pF+ypLbviwioHDm4mt2Mx+R
12LdayDadhn6hVPv2XS4s5Pt9KJh3sTqAYIFHgpk/aRa6BkYFmxmFbBBCGDUIS4XgZag0BL1HjCI
pc/kvOHXTdSULyEQamw4A0Zf0Ton5/9M4syr5bIGDS5yq7yBbmbjwR35aSlPNZrj2Msx2o/Sx4hc
YiOxV663nfoCoIB8JNdUAPxA9QXMr5dwbyZnqh6QLnIZy0nv7mw9scW0PszGaI6XQXpND0EDu7Os
54nZhh+PWaq635ncYVkN4X0y4jqRBqso/BThod1MVn5ka6joNYzYCfK5tCoZLZTyzjnhGYWDAXc9
TxnD1LynP6V9MgXMCBIvRBgC/gOtzOeCOLSgU415JWrDBUo8774mxX2j9npLdzu6aJnkuZYjzLXP
BLEZojsJyJUuPj5lZNcmF90X2TIbHBw66ULIaktI+fNLIfXXHPU82swQxusaEvrqScZCg8gbGihX
lKdkTsAIetB04slyEChQp7Hp2NEhcVMzHoIujRyioh/khnCs9RQvc+iaILABAzB3zSZ9j4oGok+k
K2vVjRHnR2papQ/sXhY71dmQEwOHRmYtMEqhsLc7AUXqrK2a+VM2PAwTaVx8Twb9gR95Icxz939h
n6Gu50BYAMNwMLBGhSJCtd5xx8ITJXBl4mw8siaisdQlRUdSXi63HumP5UgL5eHM1ppEgmUIG8eU
giTBlep7frdfQruDs70zqn7OC4FJKlN+j5ozCl/JnDRARq47NvGX2U7RABJnpIffokr+aritRV3C
whTixhSIl4KJ1Fi3Gc94S7mQ8u6KmVrSQ42daPJyyI9+A7opwYw638dF9hg+F9MkgG/R0n1sd33P
71l3dbcds8A8GQv5d/xsr9UHkb64Gro8hlMjpJ9UC23wkGBW7qVfqZdma4aU1qkhUdwFw1huEMIf
v+aSWqKrsk58Ry3Uu3Ty+fRvnrbT7NGCaNeIzztCkyGMKoL2dHiE7GkSumdafGc3HSLBmuJdxtsr
P2RYk6OjDGG3Yhd023M3JugxUDOOIl+kMzzO7eIlMZyYEITU1OuoC3/oWKFu8Q5M1WY8pOjAlRkS
77yUQlnKe1LODZMowz15SYXRL1nKqR3BghNZ3QAcEpAUSDFYgnnjWD3I3AJeMDL46zfVDOhUiip7
oawoxWjb9VFrdwsrrV1Fm6G3dNbfmOfhmjFHoAGzhh0+vlpqGJNB0nvYune8Oy4HbmR+M+9SGx9Y
hpfpiW4Z2oUtBWYIlJlVjDAkA5d5opLMsHSFmSzNR4HfhI0Yl5UE/nUEqPioApMcTVVxhILMBVkl
DstHTR+40vQD06sN3z+VpbZHdOnrP7Rn9NSKQZ+PE8KJOYSuOCharn4pqFPIriaGTcRL4+vkwGLY
01ygNrz0oZLuMz+Qq/qTKYJKeqi+oXni8dsTk0oDvCp6umxyXDWTUSNkHQQDWLNXVBfSZf/NF1aP
7MxJMLvBZ8u/rtUBihwREiUiftL0Hx9QU3/ZOi+UKo3QC79bYc1xTZ11UFzFaOe2vC6O3x1Au3o+
xqxx0kNte3HuIZXyl0mDoQuH3PP9nF3DU9HUolnLBpgFHxw61N1PfvUko2Uw1T5kr+X7BRhO2d3x
zmLetmZ7iq7FfM9gjn4C/Rte+i7/7AnrHbeKE5nrW1HVNkruU/b/9eEySdQEXc9W5R1siDTFZZz1
KiMVOOdy8nzRI7vpf+7AL1cjnfaLKtUh/yFZCz9FEyXvwPpwYMuju+a1NxNwRTMDFwgVLKfzjd6i
CiCkFjT5sHnjFPKJcg5yQqwi3tSekipKLc2gB7nWJbwEpWe828/60H4s6fUESxqDfs/8T+GO4AXB
XgbvpC+irxU11OHZdQ6cI9JkcNfss6DEaWHznJHiJFL13YID3OO1WvpGCELhkrzURt05yjB3zxaA
OFRtD0GcDMdGQJOAsuo9E8R9zrH5esLVi0vH/vt9SS9iuJDCu592ItikvktbKTwj6fT+4p8/7rVJ
tP4mWyqKimq7TucnYKU95vuZD/LrbX0/w75QudJG19OzuMQQvoEvXVTfx4ViqN2ciEycBRPbLRDV
GOCEdf7zt+1qE+Q+znEsATsqT/izGQpUIsxKrE8wXOW7s2PDr/LduvsUUIJ5ldvPRNOwpMESy1F1
eAlMoX9sUkXRMlHuXwY5D9uQ2oQXnMwLiJEsA0HSylOsNzTU3+rMlVXd/y3Zve8tKjy+JkqrZJjO
Yru7f0NyGOIoSrzFS/k8eO1aDdNqveOlm8DWL6r5qVxFMu7C2fSNolvAyvFy+Ssrxt9SSaKkElF3
FJx3Yuj1ngZd+gQDfcisemaZdrvViXxNVApZCsg4q4KLV8PCSxs8xI81Lrxeh1RKWRWt2gBooPm7
TFYgdCB09DhhWn2+TG3E6Wmv86P5bIE28fSB3AZmvtaxQI0u0TL4QiScFscl0lsES8NF7a5X+vwb
nV7ynsxq1CUfLQqvXBcEcRbd0jM17vezxRU4YFLeEmncwdCXghKBWEUizB6RXhxolRp1sK5g9y6h
HUbowzNkdFVLTlfExBW1i4oEqJ0n+DAlkMPtTaGPcX9bln6kJXlFZlLC2wTfsiI1Av1PUiYEevoo
sfbfByf6AEIWEwJcKGIKH7d/MrQz1+Qn6MLLQ0px00Dj6plGAtoRhys6YEDxtoCQiLnia2ttcnIc
STgXzwjctfM8sOYePdYm6HTY4Zp3uFxR3XvSsphk0eqrLThIxS+yu6PCdG4gyRyqRNeHMgo06ST/
SPOjYezd0IKz8t/FOHAdQmuxHR1TX86AY7dWe4vMplZT0nHVI/ki0rvWkMfib2M35zwuevHF6CI+
ngy5zgS96jHj+cUdHYpseCTn1/dha1oIKRPg9XsKR8wPxXDvNxWz5+JNH395MEJ5fYFaN79S2Rkn
3B6QMKiXxL2/enEp4Dh93SJWDoL/oX/xpxHoDGbzExWy9UunnrAZsADgYWdUxhSrfQxonDlqNDGn
yx7PAQgJmmGq7pxBQNEhO44Qas7vfDOzUoSrjCC7Lgzpxu7joa+BYlrRyFoiKnSip/57tcZyyKtl
qHpHgVzaH7LV1f3B+5yQXVepFd5qlGX5H1yEI4hd04lfIHCkKzCYAKMRv+y8EazhlAONwOutbsmj
ax+IHoapqvsMyZbJ08wrLsgX23bIpQnCPdyzrhRsWV7+ZTtVr6+7aKVhH4QDxW2aa59IribDSdp2
dPSIz6FTcUkMOLhyEG1vp1uCXTHcICLr4cx+bXNTmzOl1TprAsy9ge7tSYEnmHm+9Z27OA1SSgdw
EJOGH/STe8LN1Y7Z+yC2jC05GBUWOtSJxavzAV4037hVLG1pUbVRa11SJFdJrPEgOZ4jTfnOq3lX
pnuUcfeepD19qugVfoSMUzSGxBi2HSMPFeUYVypGTqdxeO93kedbvUddt+pN+MRfb5x7BwW437N/
+TaWHr4phdTa7vJpIIfrwwCZn8apEFcuJbOVBM5tBXUvYui893WwnYKxgCaijQHbEYko9/WHtpBa
nnQVAYeBaYJRzHt+uwakYYxfg/OozVjQyepW1ctY5bzSf8jaYkQiZHvbdSdL/eMEhZNdIUmp0r9c
+JIymtH5tz0zZwm/8lVS+Qkv26LwocsXuZqvbwRcR32M8mW0uSyrwaeLyfDUzvaSSoBTkAfM/izZ
5cesx2qxBV7NOlShHBH9QqB8wxsly5tv0fxKSEXqkrLCFGSRO3Rrs9PVDeTBh6sXCAXPTQynbG6O
EoxDo62tAQeVdVdyyYLPJCp4gMTgry3lp8uv97oFa/lKkvuoZazngIZgtN64+1l76//RiiEoKjub
lFt0DS4SLeDCyxP7AMXciZCQY0fyKI1Y7a+hkCmBoRr+h8qMtYZM/2OeIdInqQ6tigkOHkTHGP/z
sbMEPSR44HRbydtQUa0ZypXSPD5EjniW/UR/rZ1LS4QF9UFAMNU1oAlLcj41pIgIq8CL0+V5IkrM
G8wIVBL9rPgp0EQJg2yADdBQlYxlsl2IEXyGkSChEhIMxxWzZ9F4dSPmwjMFclQIGywOcIdDU1ff
FO6G6XSpCC9b8Wuwwa60xVhexlkYP1GX9UIELDFAJYU8BWRYtRAA5j01KljUssQiBPGDOQEQQ1KP
oRWT1bjs1jHW1zUjnUTdGho03pCDrP3ba6+8/kjKYejPFt3CIrQL5Qi5f96nQWhCHzTI/61Z6tPa
0qKfjlc2ECoQNenBQ1NMJIDx2i+JCchHr2N284Diw2rpyAZ+a31ixXvyad5E8g72noQcsEOkxxBN
8vXtx4lzL5uHLp3aFRNFRsZmMM0HbHBQf+XgIQROsvqgQXMYh7Hi8KhzZuo8MkHTjWzeCUGvy6FR
0CWEg2CHmoeHWozDockUc8ZRz5kchNrVgbJJ9mI44/O1PQp34cQRLEZUK9oyOthbEc9y8v+CfXL8
xYoiQGd8cvWVJ952VIi6LImydHqGaXR1FiN4PouimMQeEuCXSwtD7sfXLjaeFAIxUj3C/fCNHqOe
1ZPuAannIKNUCzLzjhBOxXvZ9cy1dpLLFqxPoTmMqCO+8zB3VITQz8cHfkcH6nssVEvHP0UAZ3Pz
cDl6oZ+jU7vnzMapZRHJvrugUDcDzMVamYD6GC2qn1W4KRatx+jygaETonRtI/w/9NgzGC/ivkOK
Qefj6d7t1xyM5w0yVkBcc0Gvn9BQ55Hw9King5V6cJqoytwCSGgHCy9jbY6j3eIcwfWBqixvxToF
amPQ/XyCRM/GMz168okcqg6gwtsw+dr5G1HYgEiQ+0zRZdHwOS2mmQYCkhRxrEKeOwHav5HN13h2
98wZWCIi3KD42eW3u+x6mjrH52gvOH2MA8NBPADsGQ1VrDBewVw2pVuWT0Dnowh2cM7qhruh9e3L
79aWDDhCjsDvfa/WMg6Bn+z5AOOHEJ4lEmRsKsIeJZxgd0rPO5jwP2/ppAOlGOYYzJ1eNFjEEfiT
r+i7I1NGvLYxAGTB7UES6l8Lyt4L+zuI9LVkTR9X4/Nc91j9Qdv/aeez10R1KUWhCQLI4T5eJH6+
s+jcH6I65/t+ZGLG/5Ztmo+LITEG2xMOuNoqq9bq4olqyRwtQAj9FFmOb8WRzZhKG4mAthy6iU9X
K/azHIss+KN9cXpWTgitlMwwhvMWz0QlI1n5Ck2tmfqrb2MQTqBIWSCzAWtNezujPA+C3PB8MRcR
vvhPIjBBvrNNLsv2JlkXP7xtbrlOvvXBC6Th1NKSsrJGx8jn1GQ7kfuhf6PawctBgo8Q79wyhfjV
AEsoVW3DEvdGZvI1Js+9PDv6/vJdT/5oVgVl1HA2rmbRqhfnxLgMMLgn/hsZ7p5m6osRqv6lrKw7
yY6ff4jqIw675bBTvKBCAWkZIVF6gv+PcagH3gc0UHBhvZphn6dDzKZ3TEXc3piirmpECGnCWNv5
ENlpz5OEsqBpIVcoe98dJn9GwZBJHmohPkc0BsBk7J5LF+KUUqdbq6Y4fogX+ZePL4HClWV63/8K
Ee4UhV9TR1Hi2imP9O3KEa7qgXb1nRZqz4ZbXOPIrHfZuA8nd0HD43u3b7LwPs5qqNS6c8iPfeCn
1sK39zIGK4s5v3EdnSwUwYMOQGG2Up8Cwp7HWUyWwU3C1XcEFwdQ5nSjLFFrK1n3mMzZw4cjCCLF
3EQMVimjAJ5PzJ83PU0w5ZwqYEfNZJ80ALXj+wdjqvK2HvuTTHJT4JHwUic78WZ8vmM7YiCh6m4R
FKfBwod812E9tpXAKmj/J8wexg8P2R3bKKG+1HqMu2KPQT60DYlS7CVMFYcsFuNZP3MEbFs9FqmA
dqtdZCdBmv8CCn/i9vZgw7dqp6vrKcrbo9qRTUUX++DLO4uK3JJidM+RL9ffNWt4pmT6Udo3zh1G
DadYlrC8UIrUDjxbfbzMtD3gQy2o2ZcjEuiZgMGTQoAYMPjhFPbi0R//LezMEtp0C9o5f5USYxv7
MPG5o+jEWiCuhb3/GAKhASVC80up+p8I0wCTH2ydqFH/1XXSU4UC/SMu9dz/Hp79Ygx5DW+aggng
sL2ykaaPi4Qs4AEjgKLEp18uRHerT2wYdg9gRUhndLtvAqpFBQWYiMmtkhSa7Cut5c2TNEo9KMYN
oBqywfPx8Rl4EGCUSYQIAGhYR82hrrcAsNrvB/+v2GfxtciltW4dsyqLl93toNd2CadO53X3cOFI
C2dnV1QbfJQTqfdy03vuSGM7qPb36HYFkx10mqO6Jg5upiF5wRLo3ca8jBAY521KdEx1RTdGekdh
YBg0E+nHexnzNW8vkTYbWVlwV4XOUQzVAmuLLHTyOncIvjEO7LIg8szyfbW7ZzXZEKDc+0L5qiZy
hTnxcLdpwV/R+CbrIFsDQWo37kbfySASa5AkB1QDQG0CZw8hIY0KUmHrhynpw7p8SwBt3/9Lg9dd
feteN8tuES4I4iv34OPOeE1kbOdx8njmgKtYCpfsR3DcxsFLBm91TXYyzaCa8CTScNE9xV/LjRZ2
RYIrYrCMgn4ozxuOoYq/nh7X1FPVI9WqIQxLQPg/h6UN3ph1eGKK7RO8GW8snC0ag5ax+OIJDrqQ
epCAKNl1FehZqDlIXxC68dz2qkeS/gZUyA7XxUaQwxNa12+E90BOECahqFbixa1AqnU+ZQimvWra
Kq5ZBCYmYxLj01YQt/selfcTweQeGDvkO0QnWrO8QQaaTlOxVlTRWie4RbJbwCHnzfEBGd9e57+t
J2swuPXa6AmMSa3rpoJbrcvdJY/gEx8HAvGrpvb220CLegDDB4yUkYFDw8aPedmlDGczU9IphguR
eCSvgnf5t3LO3SBzZq3EhfQX7sUnddk0zrgGtZOqxfVUIYPNfzT4DJuIYY5H60JNTQlUwh1jEr3b
wPkFPGnhEKdi6G9TCnYdGZN17VSTgExdJaQjkdlE3eFkrl/lso7vC92x74817SW/Ax1H7AjRZaVQ
kT/rA4ABEVQU87meL6veZ5IT1YtDUUSwjI9GcH99HSOGj5CkiO4RnkXE7IS7mxfsnYrky7q0yKnS
xRDzDF0tP+8lQQPaTC/b/iu49BnH6RJs8uLLxywuZ6VQpIiQMbt3+2cOmj9cs5Uz4gIEHLBiMBDG
vZYzVe5psahTRyo1Wuto0Ewi7lwuBFt2qW+VGfFc/X6hFzNKLb5iX7v5PX/VmDHU3Y41kLuBBtYb
eB4D6X07viBSSrZNv4oKHdgIyKHdmNE5JULsCfVNGj9cnC1fY4WTzl4v/kZJnBUA4zChyXYgMZUw
oYgKg+7683HlnXgcDndZ8x1k4W9kAf4Of7kOYvLtxaK7vwIUfuVffoOSeQBVXCQCQlAAPa8vYqmH
RmUJuuXUC+vfUY28n4oVO1MiJ2ANUfbctmvHDD/i7xOBdEbpacaRSONnPIPrqUq1ByQ2wJbQJ5jM
OWf2THvvvBVlpDzKrLTSytxseDhER/PQo/nHD/Upip3d/y947sQ2RYBv8EShktpx+QrCkqwByJB8
lm06jhwayJgw1EdLziAmxGjVsxQA0LzOPlfUGrAcyZRjU1UCCcF0urKQKLAWRCLLVGZywZFwct1D
NKeSaR5kV29aSfHtbtiFhT8FIiqIpXwnYIMwQe4U+lcEk2ov6n55HWpNvU+QBRpoXYEf/bW6m5iO
OIkoxeRodvkF9NiKc9Npefvd8VUrMMEAkyt4aYXxikayG1w8hlUu/iYEkdVjVW3L/dbIQtHkScbw
5kXls0+rehLkX2k3krJRsiOstaT92YOg4Dp2x8Qb2x/dKNOX18RYdxN6aPKyGEYz1CbIYnnUBlSo
Dh8wD+bWuYdHZhxA2JsNyMb/C6Ti7RxP8vTq8jmhTIzajfFmeQ29KEY/fPRnNedKDZ29BMXCcgRh
WBV9oUnWjC0uF3G5gmHJ0uWgQdMskbz2nCWSwGK3jSgJ8iemONpDXnLCQIWaQSgX8cWJXdhoKf7V
gNxmMp67BA/p7U/+aA3U1LQVyXVQYCaLqiPkf91JpeMt5Ub8LyjcBSzOXOKCKr2bl/hB6JhPVMhh
PaQib+Swf21La+uEAu5Z6rwsQlShxoHFz7tqNzAPc05qT3coMByXjqOHqApjki6Q2NMF6Fr3uU43
e9HuJBTA34XCZL7m6IEYuQH2GApdKfbqblSDseq1ygYLAncubuXcwHQRdBpYY/iytWfqJzZx3zEE
YlKeqp+12pIuccaAPbaiID0MHs424MHtQDArMMNmlG1pDzBmbd0QPkKF5aFEHUIHMdZPKtN9aPdx
LMZI+iAadMkl13mbLiO1WUrQCBz5vUh3rcbPCVvEauBZjhwQRVHLkbAzL++GDp/c7wOcCLc6zyjJ
SNK8j6mPvJ902M1IYzOyvtzeopVilMusnAvQd+8yEPrl8Mtq9vW44bi3cmtmYMU4ksMduNcIIfxQ
ShMWRh78b/4qNG1Kz25sOzlezt/9OpyMJHXoloFJFe2zaQEQ92vd8ZJtMF9BmqHX43t2h+M80Yck
MxcY0KRz5Sb+lAwnx/8+6BxBYsWZ5/d7Av+uC/gZruBiUyOGamj2/f/CN3xvdW6MC2wgpGk1DZ0j
JFuj7scmz7AQqmmX0bPKWInoi8I/xwoiUZzcPGUBYGsA093z9fccaq92Xle8kJZqeDLLI8aTjniq
qx5AFChS8A7ijJ1FmLNYoeBIg4VWZRL2cP6usGJrnBPDXNo1BggI3Yb/QZZGrVlhvV341WL2fZFZ
yuQKdII5jTlX67Xc0rpBtjWfCUaewVti03l+69xBL/bPR1SaK+qxagRKb1s7li45A0gETogGIkn9
p76kq00DXNKXR+FKMYJU6AfxqLFZFa1DkaPc1ZwPyMUEUlC9RkcHjxCYlH7rOYpK6nHdAgB4BNcv
I47qSPxZe8x6BHUztkI9dkn+YWLZX5r6u4cQBJiflS2BFWh9SOQ6oskbBS3Mp0uT4xTDm71kt/AU
78ZY80FP2uvnmfsTI39TiCh1tsVq5YVePYXjTYEIGMGzyzD/fdHQyLe7m0Mz9AZrJzszfSNR8VdR
+xPUFEKy5MDcO4ccwOvXIk3TBt2+4SKS3nWpG1iDL9TpxiPVnGMN+eNkccuSSZZynmdXUFIjap8G
plCErFuyZnhLpkCXcIsdfVBqRwi8sLvGTmXG2zkc50p5JUUHRRRyCtma2Gp2AkA4ZIEGjA93T1tf
XARApvN91+OcIWuvaAeaG9Zr1myJ2KXrv6A6fYnlgwFpKZuKDIn2EghidnSyCMRoOgz9MIyDWxTZ
CHFQQFZSwIWXoYLQQwyPzIOGX099ZPwZqZXiYwQXuPeU//8NdXicApEXMEcYnIifIFT7yo49SjJp
kfCwwbPoHI08AHG7bdqYeyIb4kgWN+S7xdjIjssSYb1Bc6Q6TJc6Phwkpo/N4/JXD1tJ8KiX5uSw
3UnOpc+R+5+rkFuuUs3JuCP9IPZKmfup2J0NcDwJ2l2LjroSdR7BhgDS21R+bHkZ6PwWJzmwMGdl
62v81LEWv1R88SOTJ20RiW7zU5IGrTePa4+3qzw29e6J8vN7N5z3GylhE9Q6cH7afckRH5VXdhgc
12Xif8dpF+tAqaCJmEVTiYVPXgGoG8GumxoiGaDCIXNZysc0Uykph81CF3zA06wAX58rs6e6hg2m
NgmyScb1MaL1x3iVLRbZMvQQHGKQt2Q1m8bn98eKCu7D23UHHoY7iR4IOqH7TxbJvG4zSkZo82o6
lHeqqFJKkhN8I/qgeIkoYtOry/NHcxYoafTipsQnnPsS+0Ec16DwEAv48KRxuA4TjwONg5YVerE6
HlDl+0yaya19vNtm8SKQzUattOOlAemQMcHGp6m4BjHO9xjYZtRbV7JME3XSvhUXTDxNh1GLmt2L
fcuk3tdjU8bundanocmie9c/YHGcwvLWuRxXimBqY3Cl/3grsS2WTjMh0dhpLyTDKS6fgWHwvJOf
Hduz3Nev7hY4BTlSxglDQQlfzUuSLQM4Wp3qkr93HNDuLViw2aMhhwNZy61XvhWlhDNJHg1s8Y9n
/nPBPzYOwLYSrkgsHrrBfWNrMpyDCfVusxcus/P2kWbyo81uuZv6phTPqx6iug4jmUl2H41EtF5F
XeBiMuRBAwk5NSPwV4xZ8THi4aMwrlH/fbjnQhn0MADRJYA69cduZOnallHDX8ozMZbdPisyqK3X
5OXCpytGoF1JnniDGnt5jBxnLm5BF2Sz02f+dua+maZ73E4blrbZt3OMOBmYgSz7ZqkwlcXupxKl
sGOhmptGPEwamgP99385KjvuAv09e3Bid3lz9CC3GwH2KEaB8XFqetzcbe15UivkQjvg3GemCALl
CplBnw2sO18YGJK7vAyPJTfV4lbnRzHoOP5m3/h3w3y70Mr5vlJ3fA3W++G+vEHgpKB/BeBNcvsv
CQJmfMRVjP3CjRSkUHnRmxR/2nnEbkG4corFyoNtwE+SlqItvvGjxnCOYKxS5hT1qRspZP20C8q0
MULz5fTzNzJ+jtELcxz7JEznLXSBZhUrIH40Dnll93Sn3OX+c16+8cbMtlnZyiKgmy+4oIhXxRGc
jsz6hXKEKCnN2COgdhOG/of/WGfA/UZk+JU+qZCTbH6IxjtwNUhT7lkVLdOP1HQ3rOQ9WXjLC7Ch
S/MtbfSAcOemEj381+lFqenbfD2QgRnK3dgNUppDx4bHIOzZevT85Dcb1mTtM49HUL28ZJuuG4H0
Y0N4Yvm/iQWHEvpzhxM1aWdzaoru0w5MvV9g7ljdaysYD7+a0qLPJkBlGSaZHzQxcJV/fBiK3EQe
AX+ZOGllKh+dG2gfeWkaHkvex29QqvpiAoPuXgxAnUcV4bxN1ihp1KZwZ3fLZLB6qoYubgBCVCa7
IK2sfIP/R4QuPclilKU4lq6epr1Zdu3I2NA54l0BGsASkXuQjKTbySIdRk4iR4pSIefliMkJ+xwj
uYI8NYzzb3HliHRTYqa11X1ji1WoE/hoM/jqypehYWb4QQafCVGnKH+LHQjJqKj9wuopbrKq1vsU
eqgXkr6vqWIlcVx8Oi/Gjgue/oyJiINpYqJ7N+2L0qqCDDRsRyR6uEF0qqszDl0f2sUwWy8yYf6O
WNnZcg60jPksl2D0fNUnEO7gwkOy69ZL2m3r6T+aHK2BxQex+70M2mQV2uq7RyDB5O5Oxdplt/2/
wpCaHMLZs0Ru9APSxAretU9CBSlUzTJOu4HD1PWLT/3d7dE/hVyxSEQUxvnRhrThzzj7yefcTVYo
OywPTTiVwzNUskmj8NmUsObzgyBq6/ZUXS9jv+P93FmZmccJpIIQlEILtiE4k6evBzy0fxJ8vAoK
F6WxPlhDeZbHmy5GeinIyJS7RoiDOsK93k2WMGbmS8j9dL+8DC7LnC/2lgaT4GheSWs7M2H7dL4c
nE+0U/vITqJYgxjfDL3zr0oU9ybgJEr+35xrFyABQ5ZRGw3KcRYIKAsy/W4J3odzAPBJcRV7XIxZ
uyJP7OB7hkuV7nEUjeUKNcBbYV5V1onl29WL9kdX9H+ICBz8FtxoiN1Z50gQgRtwlYI2uuJDYi/F
f6M5JfKq3+z2Un3Ck8OxDKODcGljW32/QsXwLJFjOgcFfiDqiMny7S3FUYV8Imbxcu4tBwjIMU/c
H0qGX1uvTAH0r2h6sn8r+uv50sJ48kDGENByNFY+6XnqNlvsoEnHsvQi1b5ckyCjEUjw+YgKeVF2
XQ70zBaKG2Qu/TDNlr6OM1sluPRQKvAVO7CGQUNP0Y6dl7w/P/WDQBE16l/Xwnh6aNBjU3qp9VQY
MS+99WHYsxr/2FC486l6rCdSBLqqWyqmiuXuUPIkuVciCgY6ZjOj+IogkrRQuOm9eqjck/aIBdQu
Li5XAd54E2S7qAmofV9iijgqEP50CIfsSxBOyQ97zxjNPnxBeuE55eTnuIE2MOfCZ/tTtGC7+3oE
0bYDKtcb9fn3gCLuD5QMaaMemVIyTfztsSd+NYHfIunPTIGXEx4+NhtnsR27+Kf5J3mI+h38W4rh
I/UpQzhFv9h4ho0ldBMZz/axMbfovZ99rEKtPYcT0IAnvQks5TgUhFFGXOmXCdZR4h21umm4FWs3
9stWUp6nXbU2zuldbvRMUGJeJ1C7k82AsOa7kDguAkZrLZCrRqynbBG7ycd6AQZifv2yjq4A7SW6
fMyUnCrQsuL8pwJwrgfCSocdZ2m59/pN4kk0Wy838Wwc8OFH6IqJ2Bk3iRFLhJAJ+9TThtcLfF/v
g+Euk3RJbdSx1Cuie50wLU49kOhNL0cCF180uGqCNzI/+kVpIDMtBWQd9Bk7Zb7cHj8y2PutrKhQ
hOPw+vRVt6fOeyRXF3F7ZKl9rXO/8uEkO7q+/RfTDPf2FPDNh5KDNunJfs3+90iVKAU013MMVtjg
guLuVYtoP83XcSDBm7edUIEy762foZAr5HUbLkCrJWuZifs5+/RkY0epZmAlyV+3ooKXykPxLDJA
n9MNza5ulVHw30+759Cyx05oXN7/f5j4+6wrt0YRmiIGNI2gbL3VOnxayyUqBuXF2FSiUfWtHIlk
rZnKagFasxl1DgzkhoU5FuhcKsl9t9lmhOsx9Qyq1DuBUT/hSvZh4sdrB4dzewGi6lruQxUofHr3
UZlXJMeOWjCs0Zn86gopKPkllBU+DCUYfFG3aSm3ZyWGO4uIvBAEGMmIM+yuMAEKZ9WgmuNK6Rt1
EKs10CL4pWifBfnQu4H9nhwbZJp6+Fi4i1jMPRJ/NMIFPlNEHmA+H9QMU3x+DaXXEfsNciYAzb0c
+BqdhsQ5tPXefiRTrBF/UqDSdyO/aetI6+mQWcmaNWQ/tX9YkPEQOpU6vRxqbm+njJVQHZNeMKvn
+nsw158NxJjeiqJFJa8ZIGlIAVIxPXvIruNzX4igVeGED+PdzB/5acRbqg8M7sRVJE0D7KWUY8pN
NUD/liMiVOlBgNCYolvg82mkrHXtixos+j5n4VLExcumtwv+BqPt6vqjXjKHxgbSQiwA+ZPIQjUf
v6DT7a7BVSdnPttxwhaDXYOhnLm3+H3B70xlwwA5F8T0d6YNrWnIa+e+ui8pr3L5GqOLHoOAYNwj
mIyiU8MJolM79kP6WI6ZFxlfZ8CeLSK0WP1t0NERAJFN2gl2l9KxwSTQ3VhNDnAfdennQ4F++40n
zAltq3vzXb5Hk62ZFDWxc64fuHg+gM3v0Vz2sBl+JldoYp6+0C1WxI0+uOKabQ/iC/YZPmk6tOd3
zmgWUDMrPCcnvbLltPZpllkCu0GmzK+VKgGTBSfz8AX6RYGuaOfDUE4PGPuqRK06UH3bSgVl6HdA
jDVrD9H0lQj+BmFqMk8VZrp7nuCfwpjVJA63xrqgNuf8v1kOzMJJ4IW/JpT3PyjDriocfZEcQI/H
G+UWiQOo2MuCTCcvzRPH/XXAgcIpBlWIt9RnoPxdjhhO4CYqSpflhTqiDhHbhI5kpjmS0zr4BZCj
ar9M/7oE06XHZPw16sygVQALiQ4kCS7jK09aFs43RAZzeMrSVMsnoI3mH8K/x0VxfijSDCyXTwIj
YpQdOwHny70rkWIdzxmjeEiGjnaABungPrgwXZTGsNtPPPgpM9342NAuJfYJenX2jAOQ3UKrwW+U
hiusxeZZ7ZkY2CDK1BsalOz+LlfxhEWpnSR7CUG3pcbWCvrsz7PiRFXQ0W/g2Le8zlKnQ9sYcCKO
0kXXVgXTGixpeq5YH1HUH1u8PVqKjHgqqWO1k+X+FDYndPcjyV7yXVSK7ss8iDOWlHpQUq9irOj/
O0Jibx5vbSuGnFg/tXsn3Y1XHD08gDyy+ZP1eIFd4F/2OEF28FfpyqBS04olfedEEsNDOeKYVMxr
DrHCg7Irg7DdZ/n8wEWVsUW4FqYPjrNVTWyuFG38fwGbJj39GjEsMfN4zSAI3VWXsT/tnjsbknt8
qgzsVswm5ke/1FM1OiPXtLg+zzY49oksYQuGGzG+0k3DrYRZ961dhPYuR6hZaU1CaVY0pJwl8jjL
P5k1KexrNxNQp7t/XWcFYSE8YZipS59giNznzLGU1YHQ6KyQHfjLSKSXwbk79OHz9hbLJAPRPHHn
OjsUcwW8vmCkzMzvdlPgAtfHiEYa95ZQXAcZVi/qz9qPZKGgVe+qQSQWqI3tEOvI8Oesolt8aMVr
6CkANkfai5CkdRei7vyGdpmMthjRIYkrpllkUj1tBzmo2uRLHrsYxlia2q7lWs/s5ppbfKdvO4MJ
MT8rYEUWC3jDyk6fKHFmU29ggfmgLdp7I3lvtxcF2iqkPqhIMYVQ1sDrR1QlYyYmapakSPYTqqyb
WkPz2zGBbbHBpF1qzevB9rAgDv3U3YCYZqsBduzcsq+NGj+KwGMQ0mOyKznifao9lc5FajAUs4UD
4RdE2Vh069qa5eJFbPBBI/2Y+WyGUwQ7utWsdliclAMW7UT1M17VoaMrPsHapgxVEJmQrHz+HW2V
q/G/5DUoc5ZT3gGTq3/O/Ki60wwWDH7wrb0NIpHnQl124hPZiDQ+SwbtloW0Z6vtnlmMIf43VxMg
IJpjzoC8YGtIAo0HOC8c776+JTBlp6cAPG0lyxLqQ0WxS8zLIaEhMdCXtGaHcoFshjbobw8mJS1A
zjt1fH/q/oZFeNkgD5IP4iToCDE6rHF4GrqAZFTV/clreUuuBGbORV2D7JfsIEYh2w3JHAZbnrqq
YwbdcXZUeoNhXdWj8/jrvJN72L5RC2dWUmIs/XRRtCI49lf3DMrrBUmvkmsNYc00ZfWuBBypvRhs
7WEWtIQsLQxJhaCg8Mfgm+ISg5acbIgO6D4DBmOheCpEhnLxZ7aVbQye3YyUS9rvNYKPHm/G9usm
lWHRIHA4ukRc6z2z0LPYnpRkju6m7upHjzwpHRSn0A3r4ZcjmYmh0HHrnhC962mMJBSoD/UAUHnm
YLgj6zyMsJOkglovmpKqt08weWJEk66uEFgQPgsz/Re+FOTZRQECKkp37Xn2aAqXPHnK7XHKVNKf
DN6fQL6PjFGMwTlOhUJiClvwpdNGfd1W+bbuoXCAVBVKApcLIlyQKd9Hc2shX2jyifzExS+afRSe
cmDO9yzGwkPo+qH0Rqmb6ZGh+RLeRoFN9CIBY1ok5uAHQZH6DiAykLIaSaEX1wa4LW3U8jLEDMxA
SCyxMHKW+BMr1Ho9zXjxJQSHpk5aNcdiz7va7klid6/Jn1dwppD0B1GLb8mA0MkvIq/WNktqb8Qd
xLs3lwzVBRHTi7HuwYXECN5IFICldoEv6xaT+OijOTTm9/RjSI3t387lEmqwKIwBqQNAmEaf355E
QKdhq+2ejbluXaLsj0K6LtPiKdzf8IXYDWMj0ig6sWk0w0PwepnXlcWCgETYKanm18jrti9FsQpC
dTmJxwUyEsVIeHrgTatdIi5CmYSXjQS+puAvgxZla1komPfdTjw95QESyTxnrWCcxLDyOBVDZI7l
2eh8PAUL7ZXGcvJ9kQn+QF1/PwS98ucQ61DtVA5/e2HDS+MzNl1n1JXzqnW/u8wgz+ik9ctqV+YY
2ybWfTTRTzQcwdPmK4aRZFXgeVV9sQY28Doqw9rYXllnWdQuSn/p9QEQ7hRkQMTmHGYFv8lgwM8B
IyNEe0gmnxFZ8NmlyVedpuvxqYECHayYYBhOonvxo2NkJym1HAoL2wHyj6AYw2WLEU26E3Ah7qFH
clDdjhDWtZ0rGOhJp5LQlZBRB7QgTcrSN07wJWkZAhCZOyOg7jCh5oMPKIVu9kaVJYTskw5Ak2Lm
vRIB3Ye0pDUj9lzatSyjCc8JyBwDZYBC3JIR08Zfwulzsm/5g2d3eD7vi5aCOJOHslrfYCBLXL55
aSIy5q4aaKTJtpMPUgtW89D9Uw0w8ZwzSMKimY8y58lsoZzzpd1EIkcCxPbRrhBIHPJQz+O5xLnj
1iEKDw626fT8aBanTVC3v79aXL7WiEHzTw6775dTefbmH8Jn5Y6V4nnJl7tt0LOv4E4kQ5rAcKi0
jtL0pX6FPT3ndLw4gp/0KsUw3EooKwMvsvG04n/J2L/+JFFCZOuAr2PVrWQXt4724F0Ug+k4t3yY
hbZdkmGoNm86oBcz119lq3iIxWoY4IWDEK7Nxg5x6lYM7WnDAugnypg45mMpolK493lyBjXgP0Je
mxEwktfaaQWhWSrTEcLOoC583E8kiKecpH6Lyz89nVxu+e8+BhijKu69WdrYDSH5u6yQaE8MmdGz
PJcGxt3zOAFlc6OSApsRD7g4IykvEX3Rndbiifi1ElbBXoApJCvo87Tp86clmSVK5Uy0oGMceYby
9vAXbX5vCOjzUT52zeJ1esV7uy16Lxw+hfGyrca+hsYRbMlKcsYmFWhMaqKiqxtObAfJNkSazA0i
F4C5dE39CtlDnu6sVTFFhr2p+E+WLIgB732/pZ2tY4xAmgRMxM21iwC9zP5wFcXzJZ4OM7iPT1gW
Vm1tC4sp20mzY+5D5WYJSEDdcRrTB6wub00WRC6J5OhUxHgudoQ2dnbz9NdOnuUYzvTTkF4HONGU
T7vjQLxc+bY5RtqhKEQtPgZRAMY2+01X9w85YyoFSTFvCFGhpZUrmy0XxXYE+nKEPX/BHi0XCK8n
vDkwm7iSG05ihYESqArYnj88yDyl+OF+yM3hlYZqo0Uue9hYEKjgLI5bjy45UPtY0t8f1JDcnp5k
T953vkwlFDM+Vsq4B511C+KJ5yjf1JF6N3UMKZEXMWDxsSRJxR7QNefgAWvprpCeCNWMyR4iaJ3i
8KGCGBxFgc9fBXWiROto6oI8qTf/0GFk/uETRYZrQD2iXgw3Cqtf0yB8cwOSw3ssf9eP4j5mYqb4
R4lILrz8bHc/fTcgQ6pcLQzyh3XP6H5dz5lA715AFTRP2SzqwTGfggRG5DaIIJpcH77MDCqwY9iM
RjxekC8DzjRUe4Rf5tul7JHuqS8UTERlsfIl3zhRw6nitUH/nmV3cqC2idFBOp8HFXNkRgqgQR9I
Jkp+t11arFvSdDzddP0Q6JExmTrhyWSsb1l73Y+FUdr6rloDqpcPk5NcGvOalcosomfbef92p8WQ
QO+8AltBDn4epSOtgURj94Vgq4UyAdqSYS8lz3lxcrvkdO+wxl/6OHSa/XgtOtSkP+v3As3ex+wH
F1YvN8zfUVU8kEmnIRx5v2xZ/83zU78BId5gKUTBr/G8VIQh6u5YTx5mOEYde/V06+YXyEalD6Qv
UtCJgcQDFVP19qbQwaiIWXbVmuoS50R56ps/FzCs2154jX714CRr3UmZH/+r/zFOiJa9a0HiMgoH
vWeBSDjBiMSbeczhTqbM/xJWFs8niSyVW+MHG8vF7GV0tUKH5h+SeKgomwSH4mahp4Bu/Wz/Miou
P48d/GBBLZT6oA07mJ807nVhiyZ9QFGxE7+3pPvGFGEXZmdz5sJzK1inV1WwkQyyo4FXY06LF7E+
qzQIe/ZDs+GWJ0/MCUlCFABiARcgITGbgOQ93kR6X12CROxFC0/7Y4GpucuuSJ/2M6tGMjR7hoEg
x9weVJ5mB5SLLWOJQIR68bI+gXhMLzGeU5nG/mWDYtoyhB8N2RLG8hmH70h5Z98a8gaP7v5liNWT
rTe3njYX7TXTRy+CSZTVGt4R6Oo1FBK9c5Cvi7M/Ij3PDwCu8ZUhWXIKC9FW4mEsbEKDN1tcUyRy
Mr0ad/L+oRux6oj6T/z/KEHN1nKOEEfs57kFZAkBavLNV/JULsDetbyBLZHAjIu0YXnfS9jP4mR7
VPCJ5u1ioqmsTadOxkz8Nh3ryH0RqK/6B+fnE9z32WIq7POt0rDaO+qTuMMXlpixYxo+L4vcBGph
03UvscO0tG4mI+8sZRW5PaS8zFbbbXfuAqJfsd49q8OS/aKuNrFiCBqHSvF5mmtHXZnirX4d4ym+
g1HzEdW95SWNzXx3xZnzGRi0xF1S4iKQU25h2vT1PuJ3XQcB7s1q9OW6EOVdJgrTBzgWr2nTQpd0
z/1nXW2vJeeU7639btUE6PiafBtgfyguwWxEhsT6bRuRo5sE81xEF7Oidph7uB83udfcuzK3qrCr
+bVPLYohjqjuC4Bvdq9jwcY5v9DoJjQDlh+6y2GMPrmsltpGxoPi7rSkJEddbRvKUbPDhxBvSGHb
euZI6xDIJyFPq1CJ8NjTKwRr6eMP8gLx90PLktDSlpE8Y6fDLu3ARNF26mPcswZ8hdgLJg2DkcMc
LyY0CepULoYv7b/8iyh2ZONFXbv+ty/5T+Ax9IK77urkdjm5Mm/KTQfC7ziAxgP28k5i/s9/udkR
03O82xGtFFqfAgfWcsGjKs6EIp3uhrr7OVrfWv2dSsRQRqCthTqD92IkIFYYZGPL0VgDifIBN8fl
NUszZ/tlXaHSmbsi2ap6XaNPWUM2GuZC8sv+bLPGSzKg4ken8yqEJVpqSyEeFePUH9c5FbtDRTDi
5XOUCrPONl+qVzp9glv0lsiKnNamETFJBhqwaJ3h3CMxWddcuBKyAzal0Hz2uqSDa3IXrhwnusDr
lTTq11SVLN/jTzHbEi2DMHHYC37AamabcViz8JbP6aHnqaqIVTMqplySsn7PcU4JIt1wB/fyJKI/
BJXTflqkZTsSvcUkykRv9UWAHy27ODDgU8mR4EQKhr7wU9t0qS59YcZuNVAdUX5iUUEbabKoAtZp
RwruAXSGikMETOjQA8FDCfbENnB92QfjjR1qltAv5DGopDGugriw8t3ir4KujgaYG6xAMB6hVdv3
aArhAbsmNm2fR3fgn6SeUCSTriI3Pbc7TdqbCu9vvr/71RoJO3UriR8VEiNaNzPm6FUDYuIHPAhL
W974vAV3Js6GnJ7B/8w1ZZ/gT/RuXDgmB2ZLHJUDJokju6C9/JGnOrLDF4xL5hKbkZ1RSz+JlgPI
NL0zwT2F1ThaMynn8eD2xgY5RpqCl1rck2vqMwh6MLCxmN6YqmIYQ5AdvXvvnqeVUPy04H4c2LJV
pXZ3ePllNXkQw3vWzkd+MbWINFPRwyhKy9pbKB/Df4ZCePV0f0iX02YLRoKngF3DFXv3QY9gysLF
gWuIJ9MCf8yLFSj8a6Jk4eYmHeQaeSLLc5NJgprpplCSBlztMEHhBgpujk3TNQcSe0gHCFWDlrfn
L81GUUxyf0krvLw3ptYcaW/goRX60MHXtj58uGNLi9JcbfY3GI1QAahv0Ty1sbo+rugylXcD2Mpn
pYVF+4Sfg/1C2QwbWuoRTithAj2bKs86GdGHcUzQ4ehBitGmbIGgLUNCfOs9MoeRO7oWf9gRiN1n
NdcQSY+RlcgxZs6xegZHEoN+BfV7XK6v6mSngx4hJoLenZovThhvTRUiy6lRdDvwXPTpQgXLPmXx
TJuuxA2y1+FJCDl0Vw2c6itZ4aIjqYAejFFlIK5ykXIaIqLBkTI7mKcHTob1eAFK19R95XzcXHIW
GWEJoeh88bEZLCvqMgMjc6hWS9TBsK1/SbgMGRjJtDL35/yI98RQPB7zPS0f/plAs4OVfU+1R/zi
h5AviD6AbyTA+5CYBdHKpEyjrk0tqPoJ9brc7wtetIpf629s6TzUEOIt9RoA+L2bg93wsJwgeBaN
EyeUuM8TZOCw3wfck1M44euXg9CRahwn0abC7EEAtmlPnwNPVNR1z9IShZfEO4T0izV9EkBadv2C
yV5LRwYXZJcxQXoECJIwNW2utgpdN53irwcjZvzjK4A6jjV+T1UjzQ9tHBH5+Lx5BLNhrZQks587
x+r4KiydG9GStO7QJOE0rYD+gfo0NLry7LtvH+gCmWlSE41+JftmbtDhs2PKqHol0jWr/msaONJa
Si20TOmnZKQk2O4aS6WuYBOwgxMjKnRX4gW8ulgLEH4R/tUa/6QZB/1BMrSd9rdfFK9u6LlwD5iC
8+kVKSRtYB1jQV0J+YGRUGIFRIm1u9vtUIxpOjnjUQuvSu7f2URYWDu0Za2B5vYlZjVghMT0DEmC
LrfdNKAwOud0IMSRcKF/U2rB8NPRcOZ2jVXrgnjJBZkoRgMVVS1dj4s4WxG4sr+RffQofx8gq4n0
p21iHXE2ONHNx2TBaLUS6EVLjhIhytovy3WMtohYLceS5w8wuB2Dt6Is0nAWaaAQrg4hvTU8sv+O
3Bzir4Kk0F9a0ZZ74hakvrIyZNSfLd+nkiPZDRdCR4PXj8b1iMLi427o/uMPcFYpApdvXQO8P3/2
eEPoNo90Ba9lQIId62GTL6jo2cnHg7gxBB8lz+t40Ffl5K/zaw9EGVGDq93kgcIH0Rk0fnn+23Em
YT/dijTWgJd94iDF1hfyhx7n4KMwDKXAFsj2KJXXbHdEGYS1qYwSQ9rnd/90hN2knKz/vaSKdzTy
p4g/oO4qjONeQ9iRmeOrCzj0P8EbzIMoG4WU6iq04pslcfuRyDYaQcWDIqSi0sLo1zATOqJS44wH
BgnAF2H78D/eFdDR36keZxjRAZ+O/G6oaTfNVoMR7zeAxXSQ+HDl+z+d3R/bfBFcqoVXBG6Wxs6Q
zaIbLTwUxx6dAwnLB6jiMObz697zlUEShBNzSYtD9q/jT8Zkzne7FGS4zH9o7dbkxFLnz0uaKqtA
SXdmg21CR9pxybUISLzllppEQiMle8OA7u7LXQ1iwTP4ZN2ndtT2WZ+FIOwzaW2uIBtzGAHFxTXm
9SZHFoyzYJGQLhV6BY9fn9BWbM3uj1vJ4VLLoi59p5ixqv1m4Qf/ix7xFTAaLvjjDhdd2QfwoEQ1
rljgyLDvjbL1CcIdaOZ+aAnuSiuIMqm+jlJSaqAZzHqjTz91RIaNcSHUb97SF6Zvr9L/WAgUhWbZ
Snh5VEECl/AdeUIuA99dLNGetEsNKxEYvLZi2pzAk0FVvwVZxVIkxFepmUYmmmWXImucteRs3lwR
z1v+VE4hr4ozn9Ir3hWO6giroQhUC8/PWSp01/ncWAcSNJh61BSK/LLW/jOpPNKl0RYck1ZKpBmn
PaNlCXFEA7dZq1DKOL9BLbezpo/QT2ANkMrXzxkTsjXLQIlEOjR/JH81WPxoQQSDo7bxDLLU37Aq
jJR3QoB/xOxvtWbh+ZMCD4U9sPCEgi4w8TAE4bApUthj1ZrEsNRwSb5LRHQ9W1ZdAefrYRbns9C1
GfZ6mS2iBNNAIdNxK+s4gXV9+OVgJCe6MQxHRIR1P4E7YRDzTGIl5jTyToJ0hPdQG93KYYJXiQlz
7jsaMMrjATpwLoMt4QHz9MPyi5fzI0I3IRYG3ziphHviyV2PKZgQGt7Oj1b1MJvo8hmcG9Wbog+C
4OjJ1a1vnsJyGlsI6fKp1mCLqj3lJlPeJz17JbJsibYkGF7pW1cKygWXhFokp2AJVytStortE4Pb
ziz0W6+Bvt6/OsBFl1x1PfSSdFn7u1tI1QxSgsi5//+mf5OcgtANDU1DPt0mvp1Rceo98fiHHucr
Tp5P9HCg+DLFWSoZnjCmx5Sh9zqBDsZojJ85sTPwfcv8sHN5OgywgvbJQVyiHogj9ofZVW8VS0F4
XY2BgxteHvskQEQMNl6lyHpbaXOIK+irOKsCPZyHHkEExdFhq7sQ3QAvK/YU6jpCFKuUUSyUZjyc
/T/z0XhMaHm9aWDUSe0g6PVyUfxkQ+L/2EADHexvHrOR97FSPqIYvdRewGIIcpTdHFuu4JoTPyV0
gQWTJcGh+FY6C+q0RQ7xyBJAcckyj6o0F0FcqwQ69CG6APs9lFxZYSWO2kF2bvq/o69kUyTcoJvc
wDfvflS3y73eUG9x4w4LMbaTidOXHn9rGRTcyM2pkJHuT4cQ6eRguK1ioDrmckI4pDEsJfaEI9P3
oAef08Bx3NQFEWgPOvFHCh2EgTMXuyyPyFa9TT+mHJGhCYrhfGkoB4NdAi8urx81FLm86gaqBT2b
cklaKJgU5MqYvLf0MJaikzyxMK8DeWV6AgDPX8ZWrIPzWmRkllCrFL8yyFAF4JsK8Bgbp7Hqq+up
2aGhCl5AqL1KXv6eW8sbhsEZVqICFFbCNzy8RQtPpnhPmjTjTLHSKWlKpZod5Df2301ItcDL/6ER
ymWCbK/w04PM7ZnCuU4m+ZGp1a/2SBMvBR31+tyMKCqX2wGjWKWuTxEBobC9jIP0byBE3B08vYfq
fsf1po1eKNDfilTSLEVXSA8x5OuBZY04uj/uLtTpukk0MJclefWuclu44ZRd5O0GxAdhc2o++Phu
RLRbzJxynnT9w38vPWDuTsqDMJJfR+A8AfExHT66V0ZI/x1icctyxfKaxEp8qGXw4ECIQys9LHFQ
Ks+k26oZR/r4PziL++E0TQIjx+FnKrrRoAVc6uI+iKjnPwqKTczJ6MBdNtYg1TFloXFqkWel3K9o
U88nxMcX4m6H33PA/dUihnTCT5HjpDO9y/q7VFMAYeSIGGVuLIf1WBh/ysLJDJiNE25HMq1NLeR7
h91V7hwTo8LOortwE9GNmVnroF1PuhRt+QUmwZmhFviAXOC1nlVjrTStjAyaMFbWeX5MSRxV0btT
zVq67DrifOErAi9s3eVOX742cGAXDDb8zblO465GkQcfq3HWJXoEoIZus3PSGEfFX/ojZ49yMnNF
lbeEifrRYWzsPHuAcUiSkM9DQ7Q4ps3ss+dT+ebQmBhg3D7RGGxe0QYZgvmSeqEp+5m0AryySDUM
zjnzz0tclKktE9wWD+756luAhVJYdKjxDWrlmapJsIyCEvhoBInHcK/K+nFxT8peqqtWt9Bg7g6N
HK55rEeKm9GTMjhcdn74yFu2BRd0rQlz3HmkuuVSj8d23Bn7/wzI+Olp5/IaEMMDU3lhTaE3MdqP
umJDwsla6CMK7cVBbvQ+FzDeiqbKDqGnd+PDR36cUVcX8bzDyNbBWQ9K4sSph1C9joN1zV+bqcJl
mxYkigCbLIdkTClnfTzTOzSxpMXWr2NpZYspTITdHcDbRi5GCR791JdWHaCTzgxuxETgQ6Ic7G7q
YCZH3N1JeVWRFbT74I+23IVrJ6Iu3m1DXaI16Y04XpRYIh8ZoljT7ccGpE1F/Pqpwlux7YXqujlq
wuXpDGzaqlK8vCJvoBsNYvSrvaQF45FU2Hkkv+YcgRG76b8m+40AbMlYuTV4WrS4alT8jJZWJ+wD
IRqgjlejcL/XqpfLOCrgKr57vwb+aIOXoO4Kg3r0/hW0dXCvyTPdG3+7Ktj0oK5xBpb+3QBxjiMT
IGhNsYV7Eny4rgolzLgAx/t4LDXcBXIcM0cqgP15HCtcXjAeuAdeNiAngnAhoH+rKlInDIdwfwUc
zBZMNTYYQZiYLHGEuNGfdjf9A32ryjGgmg8TRZWM1596hGZvBPCkxuGsoGM9A7PuLySFjkHNmOOv
tbeFFMTKgcrplFl2orJVAX4FR0EYE1C0Df3TrM+IWTRmsr6sE/DHF8e6IBYh9vp6hmQUmA1MdpWT
sEPWXl0Ud6mr2EK0fz7KFEufPdKLhHqVV5G/rHkkCsmz2Z+eWor4yXLRIb2m/o+nb3HpBcwksji9
G86BFj7byM8AaeDNH7SYoeuno3eay+kOB8UoEkyZTaNZBeu9onVIu7oOxHBG035KTmXXpTFKzTrN
DEDGgupKoujq1MKSrlRuwuEHvEhaA1KONjt0UpPRiQfsZYA0M27Chog/UJKbUEWlHQDBCoAVqBT7
WFgwO5IyLGHe46lCZVWjAIj0DZGf2+MlOq75qg/WtNBCJHLqQunwe4ZT9w0ofXr+oaosPgcfc13x
/AezDxEENBcF4QeggIrc8hnoM+g2mq1qR1WLsUtwUBtPyYxqGZ5Etz7sJ+UDkkozzFwTUABsNKcP
wQ+H/uG0r4IOHcs+4vrn/arX1TNZ7xQ2cfC01dHsK0/Ji1L37sdS8X+xMVhJVWZeMmwi53QDNKd5
X1Q3vF0Jb7VUUIumhYZ+c4+qJzn4Nan21qBTYdeSVdk2M7+QoctICsCfyIcYRLmZCZqnEDQ877xL
2n3npETqniDxv0FuaGXUEk5j1i5nM0CvvIJEf0mcSJMbI4PSzfoxW2qSM2OHjPtopFL3geSzQE17
5o4gZE4HaflMTNscy7LNnIt/lFHBy8B0slEqJEP2KzqQqDQfAv0OrFTuAJDOkpTcpjMosFxOpaUO
k/NiOtrchYeOiF4980LgjletMpLedqsM3vjP2urr0Vf3SHI5Pe+NfOlNHyqEXC9LTdDkJCDA3rWk
FSvtqVxoYSxLHxXt7MldihyUtGamOuvDPpTAS5rY9RbJpB1wqQEmobUDGmIPERpjht0OnmjzsWpQ
I/sAFipy79FKRtviuvF466TQPyr9hax9SClMxvLxUGJBGjIqcL/jq3oGWu2F0QemwMZTExBzq5XW
5jNKAtUg4EgTU3HLsH7cbCQeFT+54dqUsVfMqoKntb+v4RVmzubs0XT9vMCeYPuPYfg0eQf2MC26
VOIdyjGOMCc5ldaWYz1VSqF5UyXYwZ1xwwlwF3JEbwULJO7YZC0CLqTsIwdb8F3WvJsaQZVQDM4U
r7cecgudTW+aL6tGNggESEHCWPoUfP2Ko2CuLDhikmQLYfc3XB9EjecdGNe6WslBgY3nhfTF092I
4k68jaLf7BshJ0V0foWjwvSKrFpILg13UCoATItVDdcjHyHAjaFlPjk966IN22lcRyxI8iBYhpli
h8pctTCppKlIseYQy/XcS1iPO3edpNs+24ihhY/NUaPqJk3+eFuvkvCrtmJcsfOVbwWEHEBhy7Wv
ZhMbH+uSOLXnFaO/oeczyzv+qktKAvu5Wupv1GME818miW/o4SWTgXyZ46nCMty0s6grBiJlcS7r
OvfOz3CtJ0mkRRXDy35xNFzJr5fzUKANd6mhMZfvE9hH4O82OGs9QP0R3aDcCQa9Ym/EkLdHJkdd
4IrrM5kusa+fUPefucl7FfiEKZj1+RV8Inl8Y82t810elgqoH03DZP44m5ncu8+Se36FcAs26HKT
nk5mk83hNibWIGDH3DVBC85OxGQVwgLwKQF2DO7vwPp2SCqVq8VKFDU94vZF+riSYgBBCvLSB1fz
/B5xqT5VjfY+uV4/tQbSH0Uom7f6cSBe+CoPa/2TMo2mzmihpDn8XwvLtv7kSU7i8pvNLI14J5A6
uqwEVn/l5i5/yBqbo7HGZDubm0xrtHkqdGQuvZzeTI+bo662VGAXLxunBoc9hNRuQgr+iFaQc6rv
RuFA4Errm8dcY7xynyATeZivxCJPXO8FpllByyyZjIhPdY29UDzQgr44vLYo4jjz3jJ/q3VtwIS2
Bg9QNHDeFLgIrBPYQ8WN9r1GxsITcVq4c/dP8IoZ/DzkjMikpPGqAWtjIbhCPUBK1QD/Qn8pZtK5
YUnjNkNQQAs+cIM2wHeJRX8V+OtmLeF/n1AVD+CbIZUaBvSo7nnov8W+rP+m4qG/ro+KZ5SYp4Uw
bXp2IPeY8htFaXoM7BrClqRNbyBdLImSmZfwnoQrGf72fyMAGELCQHAR6YxTLglh+g9COCUuffQV
0BVRm9j8TrrbCN3pp1RkGDgAKZSMslq3IV3fOtTHt7NwsRP+rk+AiW/i2Gk4NjVSD6OzZ4mZ3N/x
/CRz4DDA62RaW22jFNJ4OkgjAksFlXL0up/LbgH09AVuG8o6WN0JnNB3J7nqO4hEk9cUvWVCjYuH
uq2Zvz+48NSq1RjAci4cFmh+ef1cHUqpZhV1YaxZWJTkRvVGpJEH99xeU0L25D8kfsWTbKyFyBPt
giQhn/J0AI1HCdsPrmdlsy68OqosfoVsmLzVwO6HEW+1d3aWZxAOgHHpAKFNbbA06eWJAZfKsumg
Zmb/muUdj/Jj+/s54dj6rN3WI9ggq2P3ypviMTS5d9J/hJupBNWVtykENwfLbgRltwxE8mtly8ep
YeYlm2FH0AZ1nUNM0IuOMH2yzAc8jqdfDCAguBTKldhFOY+YChlAQ2T4oZcbezI/aXeR/Z4MVYC6
xJix4UCNEUukDVsxaS6aoo+TBis0LXV9AANe2f07WwhAzCDMIxNoYcAfCRQj9esPwiI1UyR06crJ
DDBBPIse0HegMoozoe7W30EPdCCjVbAtTEN5eLGC8cGuCgvTulLXYEW9gopsAICK0WoToZ8NTyio
0EFZQdLKhQCfL6xeqw6GlpAMZJw3wAVfrplbyyARkxr4UUZFAJ14SWXWngUCCpk5ptFA/Qmd7KVY
n55xvmcCZhaOFOuThKJl9PVwiBRPNYHCReFKatp4gv7B7PjlrvFC5Y2D4V2Rj1rxIqmYhi1yXFZ9
kI8om+ihREEpKUFqZ/i0+cBvOJj82rdHLBCxdArDwKO4AbPbumcg1apcRllYbwyYAgb38eGWQ9S9
ctX8cYiYG0JUHpapD0zrj0/dlb6RthKh9CJT9GBpNl5FtAYkA1e8GDmDnAYH1+N7n6HtLkyXYL2V
Lwjc0hOoLL4gt1It8D6CXZXM8p0b/VAdmepeBH12qPQqasio5YHeEJ6GwiJZK6J9LtrLkAk1Hdsv
/RllXmI/D8SHO9m8TWvsPJed0w57DuV9Z8uBfr+iBSct5R60UG/THrigQ6I9ML70708FnDx+ERYs
sxWn0dXejrJ9y1JbW13bh++CtdsoKY5wejmDRqOZz29QMWg3shNRdPw7c68jxLKnjHSthdFqGOjA
tKcuv9AQ1jN8Jz1I59ZYduHKLedz0apSB1xlKbxYCpIbQNCBxM+Ag9ImsraKAkZjzIoV3XiiQYeZ
5iWSH0ASHMvWWrXKlrqSrjPoBMtBs9g3T1bUH0Eriq84cUEa7SrEZ6YNWVIdeOCXhr/9FqrWgCcn
6QxfpiaWkTfr1F4YMtutxPmc0xRkLxHx3cQNNVUr0bkA/XPeKTvWFpt1bhftd+DZhEiZaE/PHpf9
lhpu97+Pl5nyteHiyts0DI+dO0nMsVkXO/tHERSEDbzNYQSqI8+fWiYwlZ/hlwanGf3zXlo/7MtI
xb8n/vrOd3iPUDx/2y9E1qQ8KWHrZ/OzTCAd6TZgZgxAvVNrU2JQPwlcr8S5+IS0gGAGjp374JNw
2eTeRZJaCIFOSCAyr7NBaRnejtL+RpPGzLjJQvu7dZYj4oW8ihhoSp4ixKWumGLQy7Ly2VqbKmWJ
fqD0mibKWQRjaNCzgr372EP7YhvAsg8ZcNB1in21xfVigdsyIjQ0IEGW3CJ07ylFpbGzNZv7lLCM
xrCUUlVstlsxMlS9vkBA8c9dU8xbvAsdcFRy6yA3cVkwCdLUhbi56Ud04lwI7sbsC+c6emdpz03W
xWQHYvsQpIzLyUnzEi8CP6sJ1rPWZiobRcd+1RbMNxLYoIE+kxBYJWcHG5SLwbfyc3XIaRhUS0ed
gcYmi1y3KuLh8PKyrnljSzhlwn5WJh0sqvsiBRTfhx2RmG84elTTKMQbcE2KsPQmaRjZtfqYOLka
QwYeRq6BLb9FK27TuI4wrd9ZhmqP0Oy8N+jcQgt2SqK0qrBRX3mKRsKsKmkVkhRVQO67yifPZLWL
xVho3i7QviGdRz0nOq+nHnz1jSP/qwgEh6D5Gntk7S0PmaEU+6woL5X26v6HNcVuiC1+Vad4chB2
ue/jMmtL70+TYFalZu6Kan6HFGbi1xzlCVtLrktl+i4xQLG7W2EoWeuCcM66SBIrZQpeaWFezYr6
L3qzdxjY9s3lrnhlEUmDFJNA0B76kRWeknQvuFh+uHPIaVX3NBE/HMHSIiCW0NaUDOgHtGsFso1u
HFu69IkISfnlMNQal4DwEmqbfv9O7F3iyyDg6z7DDiA2rIcLUeyZxT12hHz1rr+Deq9wEjpNIGvn
CmtNvBfHlhrE0YgGg3Sp2Y6UuW4YaZ9Gk4W8pebGBJgB5x8pAXpJULkXf9w+F70TaNt+a93ydGBE
j/cQAZaaRPO0YEnVTu7R9AJsWRNdxZhEEdc6oph9CRgbHfdKIQLqJkgZ9yKx6r618Kw71nEe3tdQ
ULhnyI7uVmVR93DqKVAUTnYXLkI/8wKCCjSrsOklhAFe0/dzDdRjVynQWxAAHq1zrMapneZXRmY1
LDBFJ/TJt2qeaV9KJMxw34uMrroh/RwNS/hGZ4Ld3vjv99PAch6MpO2DwEqlJpmUedNh+Qe+3SpI
e1QahBu4nnMCgzjRA8KtIX7MrE2Ts+Qaw+WucwZ0dnaBT1rg8xW3+TK2vXKRYiAFrVEyaA+JtYJh
qMY2ifcWyQ7/EbDxs0ZPhaq6BRU/j0XEZjUUjYkwxa163sjU+MPX2b3GjmOyXVxUlkr+4KWaZVvN
SRGfvtWPjeDkkw0b6mDQEY3N+Z/BsyrzmS/CykHw19HbM0lTp/tTlhVEs4jDCOhzdJoWtDRqDEmO
4o4OpM6KQ1EbCOdurW1AOqrqCz9Cj3G1IDBT8h+x9v/7SKh9k3pFpZIIB5WOCoNTHWLOnAyow4hH
0vjvjhblUnoK0tf3fAsnAYsluKCG8WVtkwTNaSHqNPDbeZJ7hYvyadWt8s3qoL9IY1QKB9UyzxxW
fQKB3Dl+9ZFZLRHE+FYizoJzvw9JH7yRpKmrarzA2L7w25wmN7vdJnlBEVo1vJVQdK7pxM+F/Fct
9dNj0XjwoY1JbqTVfcV3+tFXvyhO9ngpkw04R3tCo0/MmitNIRkqV03R6DXzTyhOzDPDKfGmvAMc
VW6biGD/KwuGEyaFjZwcOFoUbVL5JpjR8LAAkae9rScV6QKdqOHdHoS1nDSUNQ2qPTZtPWgq/WlP
fmLMIYSBxYv+gY1/QVxqIcJNVa69Bwu7Qgdp2tCV5fcGM1QxjccfL0+HmRARNJJ5JO23rDEYS2rI
oNJuoqlfzDhHS9yNPubkD55G8ExHTFbpELNGBcKWuYtRhqG8qM1wEJ7L/4Nwkoyx8f/52sy10U8A
/EsbLZ0L2lT+OlaGz/0UZfjZ2EHCy83LVCiMZmC0WqJYbvhDJSK/t0rPcELo889HQZFrGOu3XZVi
WFbEos4ms36Xg4sp/cwNwp/KkIoG3lf0BRHrSSdCGwwowiTj026sgMpZBPdF8yxjvjQQpBsecEh7
12rOa/PPw8OWkO8ghfjozfu2j4lLl7XBnjXuxNHOaloYiLRRnMOzyywped6BNDf2h6YK6KjJms6g
WaTERo6B4YXZnnUuyMIVkYHsxJJ8TAazu5QI/JKPcfk2TSjpwpUnODql3fn/diybQknj5ic8hoHP
30ggvfC7xB77KgzomFyVffwR+G6JwC6ZyIkWmqKuUuoRYkawRhnQmKXTqjU7hmrxfMGbVsWsWPJK
ZhaB0GLAF8sRKLaYl7azIYlBZ13qs9olh/LQA/Cqw3Jlm9BZ0H6EKKwGjJEbuBhnI58XAyXtSS7w
Lr4iJ/5zX4L7fAvSbtsQKUiVXyXGFHvHvawxdXOfICwUTizBAXqs6/V/bnTeeBC2+m9oTCXtcIR7
1Xuofaq/MTbehEAzIF+oNd/hngdu+eobA0tlIJGVscRbLrV6QvTvJiSUKMhg/wVSf3mF5w5l0Ji+
QG2h8ss3Hjdc/Mjqgq5+tTULSWpkJxC8MxAEo8ouPNld8yX4t40vbwQfdUhQIPqWKdIHiPV0Ib9y
bq5DvWk9JH/jQopQXEUMFWaEeXAwwSUUrqXtlBR8A8dyALHQUacMdcTQlUPPOBEg/GKPR4QCiZZ6
EliM5bnemOD4NYg3s9i7TQpamgEGaTXO3lLSyByvQXpYV4psKRuEjAP6yTKNVq4nbgWvxweCisrR
5BB3u5er7/t6PS7QErcZcoKLcCv/3mCTM0eLNgqlbxJFx6lS/iL+gkr6QrdvbZYgr1uVt9mYMsi5
fVD2qx09+ngEPD1BEl36YPvXl68LxnEt5ZIUb5MlnJQt7L8EVwoM0AlzT5S/X9PmS2K2soyeta/q
Yw6Zc8XkjM6TV6HwffPpBBnaZ4bRQKjjyrA3KlD/Tc9RBE/F1u1BVEU5tC/0JJCHtOdtimTau2Jp
rhPdLvq4Qf+cYTR2/Eas+Um5RLPao+PxGOPkXjle3lo7HoYiw1CE9/O5k3S4NCxfECFqNqoUyCyW
qUFwprSdCwkeYXU7YPVrjkjo7lu417McTzyqzKbq0gWhuXwK2iOc3zokfh3+xjFzkqkmh8SFLf2P
0xHrj1plbEquJADzw6YC/6+REyh0AIdbMnWDKJ+NhIz8C5NOXXSLrLBNpPEMaNuP1UhVyk8Sk6d+
J2alUwtqE2MN8ulhGWGHbUH1yvGCQsXE+fnWxP57YrNt3oX0MoFSDCXLWK2MbRDcAxSbApg67ydS
jF6EhRMfGoJVtRvoAQ4DtZ9tgoBmoJbvfi8dsbzl0w/JuaO2QXNiTe8J5xEP69OXLvoshCiwmD7a
3S68ixnAW/HXIFcOKGsUDUgTY/PG/FrIFu1x0SPjnmaJMK8HUEuAxgjBv0aYFXCqn0EZ7FkAuWpS
bRrV0u79csuh3tRSkoVACKPm2c0CwGg0Zx9jjzUn17U5eEvDeljtbMIAyRb4712jN0wjB8KXYrAq
uhLI77fEAUjTgAHHfdIY5i4rhDcLUd0gNe7dnBw3vW7f1aOvqvJNM2qfaaaY9s3/PXYKDKk9uscE
Yojn9j+G8XmFi2aYK4pPKfoz2C30VqdbadH8EN9gyLQEVsfhK86gRplp+19jPjnZOhRtwyuoTP/H
fh1j7xf6Jo0eEbxxMDBtqJWe/CTaeJ/bdQARq6Hs1vUgXuDLp5Je+8mRxriiddxizBSA2mMdpwZa
VbVLdPN6CJDsTeahq1kwQjzayyEa5U4blzYhTIzMShUEsMXRHB8bDUq5h0RbARslV9TvsfLKgOao
wxmLCacmwUtkRM6P+ctqpdJB6niWqaoCRjueTBhlWdAtNZeiS34eicmn6dE47sI2wUrPU6FvWhy4
SHLBabvn6e+c/KGDof9nvAgLwD21TgatfLGxMAl8XjQoOMUm1vSBFRMcnLuDLioQEAdVU7zeN898
pambrOmj3U5dCPei19qo93Yc24USNxD49HHDdUmV6c5GYZqTE6vbTjgQsthKfzvwpW39rLncf1xq
sVjJw5+QBWFP3GlHxhrGziO5Dwxl+/HfMaxP0wmNmY0OayK2UBNhH4SWkxBoW+wKECFRbpjpSiyw
op5dUsjGFWo+beq+QW+kp7MCYP/+RhKDdS0jl33V5grbFYZw6S3f1M8CUnDzHEgSkLe8n0xgqinW
y/TNYR+w9ckMJXCMX52f/3kB/tXHUP9i0c6GPBuT5IRU7cDAYhqYY4PNjZyS4BH3m1WldUIXu5T9
5G8rzelL6CzK5cbbAKa3JV4ZzfT82rPDL8HcjirjItuN7P8XWQs/kv+/sMgTiWK+/VF8HnsEo1JK
aTpb9XYngmd/4r7+iksQI/kV9XQR7tjBpf3fsf8rq0PuVDJ139r8c4uJbe1iZsMNFcloGHKx4rxO
1ZRca04aAMq6UPH7KN1KieI9LBdVDoJYPZD4RfFFO77o9JkS8tzDiC+j45HQlvCSDsDqqO6InjdZ
NBwWUSDttb3Hs7q7YYM2C0AZ9XqcM1bwFHR95YSEi0B+/aQLJSnejrp4UCZfJURgbWXN5dtm+Ijg
CdbqReC8eo9w/5A9Rk4IX+hJe/QdpSOQPGWDNJUVFN772o5qmqC0mKE8/yz7Z+JuZlqv/tazyyKU
I/laXqjj+KRoRhc4CHDSmi1j5YljiXSBKUWUs6dhPlDfEZmEhgvOf/MyBqzbf0Im4rQnh4U3BXXJ
pwZU+SgP19PYZOfX9qLor5Iw3b3hS6LyWhMfki+JfnLBvJrzqf4TBVT6fbW6vhhitzJwKmZ2kwrD
ttaLtiY5MDak4HZj75qWipvyEl83+VhHENaTrS0GtC7Q/cwlvYOU22cUOzb9M45q687JxsrmpEmw
QnFhwagUZZZ9O+iOQOyoD4tGTeKaDpkZJtoUjjDnKeIfvKKMMl7nBUErZ7UAnMWYkF/cIKvww9Sh
1+HkWtvVeKDvDoZELkowGbWAoNTI7Jfkjh0063Mt+OZjBqEm/0oUjr7UYssX9bRzTTEDwVTy72B1
iAw7/+WWrg+8lmujsPbWvhkop3px05pGwBB0xPnjRcEQaOC6XFqvNijaP3/ihaD7TYPaZXD9yyIo
voWXH2zVQ+1w6Qr21kxeREf6Phgxj/r+dBmL4MEo4V+eDNe65HKKq5/w/RXcdPyJ2uqIN1uQ2pbm
lIgxU2o8Qb8EtLofL/AvEY/kAEWTCt1KKJy+vPrhTY0EhWBdtIn+ZXW2Zg97xuKfMx6tBBNkLqt0
eHOeoAxBfCiPrz2tuNL50onMuoOmMVdRA/oi1WiD7vN7vd9bAUC3UPHXwpjQ8I8Ika7Q7Qtf6UfG
u1+Kj5qAXRPOiwbEAtavVe0jZsIkpT14n/Gq81xYOy8PFK8ggoyOeij3Zyul73cjNg5hoigm9pml
hQZ2mBoQgh/a6Q9r6EhdMNNPDEZdpI2TKmp+guA50xxPlamtB8ImjvKHUu09KobuAgtv/gLI5uqY
QK7v/nXoRHtsOUcLeivSz4HR+4PS9q5lj23bXegvTRqUZHWvcFrAT1z1y64mPLKr19sRVJoX/SmT
yJI1RIEA9ZJSFmShCnZOP9y0SuyB8Ku/6ldN+IgHHYVPlNg7yNzo0Lhy9f6zyD1xL1VZN1tD8rGL
hXcIFHiZxn4lIEBL37BXwv9vVzARgsZS4PIQ1Sl9GWn4hTRuU/cpEAo1MtVLX98BqIsAk7DC+LD5
80/oZVwm0Fg+hq/rnHZM2lGJOpVeYASiEyzKvb/+6W9Rq1x2VgCJlbO23ZrtuT5VyFXJEqv2MD0M
+1feLadTWdZMEvzKpGXOqE3bHwI0fOtUIg5cpkOljhVRo/J3GRPSNzDUDNRuGJZmNOVeRYwvEOX4
fGkWb2IZaash5j0US3lvi63ALxSo/KZ+GS6rG6mWl4P/RKUNBS2cHhVe4/gX7NVnSLg5iU9JxHQz
MotoULWdhHS3rCIv1xXG6KuYCZjdAyTuzAUGid96AK7R5h62AtPwinJd0eXy/qxVpLPBeylf68Jj
ejZITwSluDQeY+W+DY02ZR6ks77WWIv1/fLT0xZcS83WMB1kLXmHqpKA9/8cNoDWDayY0272TfAW
y4VgiCPHVTqSKSnIdWgXhRVxe9S+VqmU4VJZxxka4CeEwsI4c5AVBQJJv0u2uFQSucL/KulIg84v
z0ae1SO5/ZrqKc4G+IC8N3yld3nWbs/hkzeW/bfMLSrlSX5GLL3SOe0YXld1ydyaKAaMBB1YWDtt
8kRQ/8ogEEHUjwmSiA/cU5u20509uWi0ZcSbVqFtI3ezt7KREm4GxTeADw3Sksklw34EuhtHmI7r
m7+hxY1jFSICyscNmcwWuc/izuHzGR/MoJcZRCDb+lsYHUMjyTznenOuT8ZcPYr1kCl6L/TFtOvw
BzGNAF77RzyL3NPydD/e6yUj/XSjGFivyP4HbG+fcDeaqoDNmQwlAZYGhLKaisMQAVuOCC/12l8i
NjLlIl4Qzj7E15hFZYzuF3hIZHlR2t7kK0Tlg2H1MmWctAJGwMY4xgQCqqqXb35D/ujclinC2WFU
7V6j16oevRK7+oWsml/Sq1OTYr/WMbtHRRydaz2rPhN0dKIyr0iixDja1fn4iV8PdUnoqEsLfUKr
WIG9g2dj58B9Fsansd/UwJVjMp7UL1XMF//O174N3G1abnsDbK0Eh5/hEs7ZCDJ4VIftDmdtplpb
EMSD1ulkr+2RsTzVpeYUFEh8I+IuGfel8dnpm/3RxD/ctdA8gn/VAq3ORtzxpekXo20f5Xy0AbyG
32js4CJhQKS6dCLhnfjmJ9p0IVnalpgTnIlWTqah2HAdfiecqDAD75SHKGp+Bobd7UYfdZxbeqLI
A3N6UFSufCm1c596j5M0jAQWLkkBin3hvLGIGzOsCnxIFN0GVu9hHZ7jdjLfKux08pUmeSfk8TlX
HscgAOhcsqkO90lol9yxtez19SDin825eEaejLMywNovn5bHNa+KTG/6ftpO0pe7MpXXQwahVyz7
i7RoxtGEpwqoOIZlpC92knMmYa0B83hbk6/HzckWa6W0ixuHYoHs5N9tmck00XjdjGUwK2pfdVlq
bXjWFQ0eSRWXCiRfPw4KWELcSVzjfbja/tUJn5kFsLsTJmJU4GMnMKhRFlBImXUG/zKzriJAUIIb
gcUoyRBVbgnhpPUvG5pwwE2sw0B6fzVxWJ9WqbB1hxHyMIhDh+O//jqg9LmTr9etlPC3MiWjYiXT
j0fpS0EWT5GxgVDmCYBjVQalQqYwKPKSO0nvxnsp+HkEBm9rqcNJqMnobzhAYMaSzdOKKVqOCrpd
un+Fhgh69NPi97cC75f50VkCOTz1FAqtbAVDmA5331xmRZXBV6ENBffM+PjkKxDEH272tMDBohTV
7q7ojbbELDJx5XoxcCJCgYpLUnuiZiARzwSwnVvjwLsMPPvb5IN5N/YyOHS5oMNxh56a6/PV5yNe
IY4c8qKaoFSelCBrH1O30amGqikM12Qz37Jl7ncDO5qG5oO+NqP3SUzSEbMTc26wDkTMqVe7tCas
3Lm0TAJ7+YwuBwWQEIYM2R16Cdfa4nNvqIcxLAGjTFGQSVZtC3o9chn09gA22KEt
`protect end_protected
