��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����E�"Eq��� ���[rV#��d��S���8�v�8�Y1u|�[��_��(�\<0Ef�,�i�����S��o~�ߑ���Av?.Wx�;�g��D�����.6F{�uLM�yw���6�E�0����u�\d�;�;7M�]��ʌ����µr��*�*��Zw�)����}5�(]���>�H�pѻ#�}Dd��DE�����r��V���b�ݦ��#���N�U�~	�,