��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�I��9���:����wKϾseo@�
��5�8J�s�˨!x��3�yt�O���(�'8���C��O�y�ӏ��6��G�6X�5�
+�����E�$
�w����j���ld�$��p��?+��&���G~dR���V2�R�x��Z�&�4��a/���!]:�¨=��馆�vy�z�=v����{%�����a�#�,Û�RF���J��B�+wǦ@wݧ/�\��X]�ZY�K65T`��X�Ϗ[�Kj3!A��,ƽ �J��F���I3(���\�5��[�[�(c��Ukd�>P��c^'`	�Ӣ,��V�쪴��
�����ɢ���m{���nk��
���ʧ�m��+ȋ���,��E�8�L� �f��#�K�ܢ���Ob-dx�8/�hR��z�y�a���P���g���/�i,������a�l���O�p9����A*�����3ſ�x�`�B �#�
Z���!���c��J��qkɤ�;�J[x�P^���S��
dۇz`a�����dI��O�N8p��Bz0O��z�2�B��t����?vC��O�/ w�'��+��|?��(j{�:
��0�AD�w{8�q��A� I_��,R�aP;��r��ׇTNBtǼYgR��nHq�Y���a�ݹ�� ���-�r� ݾ��1J�W�FJg���t�aJ �r�2��jT@�9Zs"���yWW��Q ћ<:=������X���T_I�|�	� /���/ ��dd\���L9�\$�yL5�j��t�"Ȅ��}�]f�!z�l����Ī<Z��8>������0��w��X�Y�T��nʞ8o#�ߖj��ŵ�1+��Q����9P��pBXo�"�)S��\ݕ��e�L��'�w.�wC�:>�����%��[��C��z�
2�ُ�,0֩�3j�^��S����ͪ���\mT�����^_������.
��ЎNW�(�$~13F����r��� hW������A�UR������%�gV�+t�M�jc�v�*A�u�4q$���8Y��}v�i��z!�J;���v�C���B�d\z/����|���]Sۦ�'~�T�I����
B2��s��^q̓�(�ߜ��[-�p� -O�����Ǚnٸ�?��[Ѽ�@�u���ѱ�x����@Eg�nM�h6R+ �k8�V��`5[է�|T����d,l��g��*	���ԁ���Z�%��q�0��H+�h)x�斪s�[��0%�]�:D��` �)H� ,�i7�}1�O�V+j0` ���Y�)V�q����)�Hmn�|g>���آLtXVa�^�qT�m���c�AV��ި�B ��̮g͓�nZ�	m����hS�k��@A�QV�+�c�Ƞ�!�/�P�ʹh k��b�I��;�������$z�}��έ�W�Q���J��g8���9x���޼C�%�lϙ턼�&��\@G 2@xP`Yx4�~�wR���wtXX����p�G�&���k�%"R�V���&���G�������æ��|�h��ֻ���l�V��� +�J9�Mh"���pM�L���6N3���޹T�������W�
66%�#w���C�sJ��X��{v*�5�K�C�+R)? �^Z;�
�}���Q���'��=:��`����k��:�Ō�+_6�&W_S�ŏU�ڞ�o{�y���2(ʟ�JD#*"Vؘ�#�u��z��9U;�?FM����Xj�R�_�h~�$��'^����Ĵ�K��<��#�f4��g �s�}��n���G���~Jj[�K ǩt9��	��n�͵L�ߜ;AM5!s�c��ʛ˱XJ�V���q}�D��fv�GB���g��R,�T�ؓ(�aA�̩��B�
o�e������(
����w��*�Tl�bT������M��� ��wA�s�"S��!D�Qb*6Ґ6f���yK�*)�B��B;׭e�ޟ�/$�X��, ů`�lc?�
aN���=󹻭�-j}�)�=C�����$U�Y=}�aG �k�H&�i O��Gi�T����u�{��b�/mHW�~��UL��ݼ�Jx`�`I7�0�nOd4"(꼍ٵ�zf�� �m�d�Fn�/d��\l��5�xEw���c/���t�pIԫ5Oͅ\4�M�Ox��P(fִ�E�$�S�-&)����d� ����cO��Ou�]���A���}��ne��1��w`��U���(_�~{]g�1G�Z�-��_����C&�fm�\����H�C�=�;���,�Z�"�)?Z$�S�KQ��"�*����|h*�qH��ND7�E�,�w�g$���;@�7g��/�=i6lŶ<��}���elը��y�9)k*�.���YۘN�����n^�M�sjiy]��Bb�Nl�߸[ǻÞ��M��"lS.�����X�����2�������Ph�n�4sP�g�tt�V�(f�di����I�q"��D�����M��G���idF�7�3sR�(P,b�ᆝ�%O��cDr�8�G�'�k�hd��E��2N�l�1E3��6qʨ����->��7��\t%e�6Q��3l7��#��cs����ҝbx@��R���?�����A���D�0��$����t����cŁ���>�8\���u����x�n�ua������
[�S�T��6=�:���: YzLE���PjV ��Yc	V��J��CM�G�&%Z/������;&B7!�n_������Dپm{o�Hc��j��Z�.���qj,EJ�Bo��Ϭ�P%5&�&U�������Dit[f��y�B9�:p��V�%<kS����_ �X�C�r��3�;դp���7ز���c׼Ś!�G�:�����T�[�Lws2�o���G)�m�<_�����|i�~F\$���������vkn6S�ru���j\��x�J E���C�9<"7�۞����QEs�\U��J\���	�X^��SN>_��es��4��MҸ�)n�u&��67��?qc����IE���
}�G{�Ǻ�ꚤS��p�-������@h_��jSW��Zb����ף�����%�t1��#|T�Zj�v�Ko4�>p9��?�ȿI���Vi[�J/E�ސ���b[�Q����cc��� �ou������9��5���{_��0�H��M�u|��;��|�pn ��?��Y(����=�x��d��m_	=�:�+"���ɩ�{l�p^���o ��|�>C��G#V�S7�+SL2�Tg�S�m�9I��+�ijU�G�KzmT-��to8>�#��6fj��ߝ\z�Ү�3\ԓ.��&4��|�i��.'�M(jd=�H[��C[�#7���Z�#�O.�6-�_RL���ҝ�J��ѣ"��.?xW���	����y�9Eq~�h=�ã�~�珗;�~���J�b��[|4������!�����Xm0�F��͇���H 3�ԯt��#m���xi��ì��l���ey޺'�_@Ri� ~EC ��)Cs��Ȉ�α�4�j������P�u�\	�6��<�ш��@"��J�ۜn�-���,ᮜ=X �*)�����8�~�������jm��B��4�I;���ʨ.�S�F�ެi���^�����/��6�\�i� S����.��dCtXȪ��7��<=��Jy�a��C;�٠!5��.�|=#�~@c����I0͜�I�Vu����4�3w��O�@��iX|G݀�ӥW	l�zUTɬ��:i��A�U�&烧S�+l��&5@=�����!��3��w%|7� ��cm��n�"8Zx6k ��%�W����}�BًB�`]��I�X1���$�Г��!JX�m� �y�4����ba��k�\�8�7�i�ڃ���q�1��zR1|3��͞���{Lӯ�Z��l��^�x���V�����9*�}C�"��`e͈M�RYB�6�;�E�][$V@}Г5��.���]���haj����e�⻵3�^sr4���R\ɋ�a5[:��#	֣��L�(�f��:�7���E#Ě]�!_�Z�
����׽x��>����}I�~: g����l�c(a��ǲ�� ����.�_i�q�#O�40���jRq��:����
��`���]�j�k��ڹ*3�=fè,&�U��[~o����i�]�!2P!��j?��lPa�A+㈋~k$RB�&�^���<^�g�1��w�H$|r��CSW\�k�E��rP�6ӹ�Ҽ\k��(�_`��R�W/�	���적��5o�<}�[�m%"Ug��w�i��1��&�����3��ݠ��A�г~P�1/��i��������.O��5���tV�2WC�k3X�6��Χ�埅&��9�o�V��ֶ�!�g��	5��~- x`�f�ZJл~Hw�}�>	IQwq+U�3�(�Iy[�����r�Fi�Ƣ�H&����Ѳ���bh����D�n�t|��X<��J	��6��UZh�_Y)K�������ق��ND �%AM_4%*2�l�S��+����g���=Kzϥ͕��v�W6�=L�ʞB�B���p��3�f%�,�/'�:�A.
M>���#q�RI��FV?=/A�,��H�4�����Z� ��[�X�l�h&�(&d���_�h<6�o;�s�c�!a������L����Ԃ Z�G;�g�@��e3�^i��g$ˠ��\��y���	~���m-a?�ޟI�r���UO^oG��߳j'4�� �*W��W��|d�C7$�B.UH�H�Ҫ
�q&i����@�.�g����pT�	���|���k')lg0��f�|FE<K@�?.�'`�/"�Sء&OT9��ŗ�Z`Q ������o�庉$�C���!Yn�����x�S����q����&�;�D�w�r�@�O��81b�O�/��ĵ1�a>s�vo�,�$�<V��R`}��A����W�Nff����VU�z�f�/���EFl�^�J�c�3���6�J���VK3-CkF'�@VYY��+0��|��z���o,��c�'9~p��d��"E��TU9�lf��${�����N�T���ǣő�t��J��~�*�����6��jּ寇Ӌ���bA��E�^c��