-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eCuTf7mV7o3tq4my83zh7rfR2lI6AFwtxVh8JpY443XvYqVNVBe6IqUVlXmG/qIuRmcyCJAwsIHx
oYgnExVyjibq3DpZ8T7TkGOq/XmxsOpSNXx61PMSODuB6SGMbtIQJf3VUAvtjW5Nfd71hRrfE/IR
/Y9p2uozpKwRFjEavvy1fbPXJDii3ycQlUlc9oc2aWpOLlAtveHkFPfgws6sL9N5UhsLvyZFb5Ou
osANflFVrlmuGKm4wE80f147fWGz+dnFOhGGNM/4yOyywvSmpDP1D7RsIsqe1233TwUIH1rI/gR7
bxuFsvN/Y550iWU/Kdc8Hd4lV+Dcz+TF9w9ArA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3616)
`protect data_block
p8Fm060+Z7AAPTuKVZyK3FktcjFPNkjh+vuGlS0ctp5Q/diqGGehqAp3GV4NYS+VSe/N4zOFe/EZ
xmvrs08klq6w2KKUOaRPLRheRYgoM+iTtctwkrF3b8AGEFFwBq7LF+W2LTIDDIQoCMY/lwSIUloV
u38aXzN3z+Tx/z07ciFbSKkl2TeKlcVfrSzBE6G+fKSm9FBUKCCih8GC8LtlfJMPgo/qKTJz88pY
0xpwnpXFYOviN0LqUAzlg4JYJv5HgvwuJAxEfORwr2KJMkIWq9gxD8hxbG5ZVwB/mu2IdeooEeD2
YCEqmk9fmJtHxUaErbqWSKnbdZGcCdFy/SRuprsJub6j5Jlw+X9v1e2bEWKcguoGbowJjoB8/742
K94+Ltp/GWnuLSnCuVmmswbaJIa0CpmI2/fQtUtznd3cPLT2WjXy9TXAuVlQZNLFkQsXCeYb0XDs
+yOJQ1FvXyKYr6SH/ivPK+AbEiD+xJseFqkREZMtNPGjtsR2Kzbvwr3qR+JVmWhah/9fT/RHBMbh
+o4QCxr790o452yxc2DaQBhDVNceKuob+fs3Om6Gzvb+DfoSZV6xJpLGGhNZvy7gVL+W8Mda6V37
4rfFwHb8vcHcuvt4wv1bdOdaPCh0sY2eWZKsPQOxcw6WE7xBnRwjX6ZEvUE9JZNQLw0DyMJcfOoN
Lym+4xn2OalWrpk/qdEbtIfrV8467aEQvCT5e+5mgi0rOV+hezC4nfg/ZL/FZOESHmnXgUasbPVf
zGbuHWFANqqY8ZEOq/zINR/R2vwb+YivEOe8yNCbI8NRdRCbURjRGUUagSAp0ZVG5/5GS13/A8wr
0aqfKwtsEniWFaL/61YGjNfvKwj6V93+ax+vHjMFk4milj8d78eV7FeSrcfGw8MTTbX2nxxOclev
Jydt6hP+Ypvbw9eduejpihxh4ppCW9chyc09KGsbmIZ8PyVsXwq2BgU+4zFuVC8d26kUoJs5hHp4
QorMXoER5oxaD72XLQN4XO5GaoMiLluQPTLN+F1NBpsJZM8OaGmZzkIInhlLdOPaQeV9ly0xW9hu
4pP7gZCz9i6+ipqNMRUg2mFZKkpbES0RjU3PDkIjjJZ3g+V33z+O4SI2Qz3nrB1MMtxVMYmPcu67
c7/prFXmRSHJHUkfQlnYsWvJdCwONz9Ccnhl6V+xYhRzxY4KHpRm8bUOlzqVpp362kRh6Bc5asaR
1x1NvqLmtphnnkY/9vQtA4tTMSfujV7Uo9XtsuM1O6KJWcG6bf6Ck+CIvgHAXrf2c95IJ45lrvcB
hdr8WT6/Y6MJC4q1+6UrJn76PAass7BdXDj6sgnWnSTQ1k2MWLvnHCVKLNwf63PpBcrAyeg8VauF
zwTVNF1nKT2DKvgQPzzK/8mbW5QYyMCurSSBjJ72IKfMsiu4tUBzi8sJosS2RG+4syjfLzIQhyrq
ulykZyhRQQQRDSrIPbj/HAUmp3o/rOI20iP0g+/H3TRqRUKnK64zCe3YkfyYVqDrsuGBADNkinT2
y95FXUGZoT44DjB2dkbmdguTBm7S0M6Q7PdOdtEA+rpcMLfz+D0/Muw6hlg7ybCdcwkREd+mYzET
sAfsaXkXR0yQ7GypfIxYYexzXnF83oDI4grVL6mSXxcx691y6r2MV1SQoN9vP9kHey2u1wDKpqBH
AZJSlqJjahEvaHHGZVkU41ujN4S1FLED2aP8OO27Bj6hNHpPGg8JWn4Jht5LvatZ+ze8d5cM8vqs
hBdO7Y2JWnPfnp5CMr0WJ8TlejC2mErUB6YXtvGMoWwY+7mnbxymE5FTcsapTmdnGbdfp7CX2Lq4
K6huyqS2aeyjjsypWYYj6A+U44wElkIVYxiHuY3YdmDeHZPhaSaRtTs8nIscznwVmdms2z7FaFAT
7l5CcwU+I273oGKPeC7UgwE2tq41/PQ3D0ZyLYL03zr0lWQxJzKOz5W2i7vECXINwh3Ntu0dfSUI
NXQor+h2BHWnf+k0ro+ewj9jJOjeRCGMYSVSmMMXnw+uFeJr5KgsW3bTWdWMLnlULUi6EN6ZgWtn
ysaBUbJ1kroqil6Mt1QIzTq/vEFPmJApLJi9Mk1GlM0rUU14yrZgmATi/AdJ1WWvur6jgXCJRly1
fB9S8rugfuIkraACmmG9X5khj2OoEp6kMPW1PpoJCceeZ4KVSG049hMnMFMvWPn7r4RTkymKK4HS
b74bJWwRlfqUW7sBziBcic/gsuizNy/6zVdFgsInvzWdxloMuYBBPU7so6IO7fC/RYKsBtPxYoRL
1ktCw/IpfheqYm4lW7rwRrSaMZMPGivNE99T2g2cIOFLDhpYsET4cvoza4kVPsYT4sUkfesWZhRa
NQQRndaV9esYCuXlr18IG7aTDj2zsFmo3RlHC28/XiHqqGifXsdSKmXYc9VA+2gtu2gKj+6bvia7
3vdV4NQ8ZWS2jLTs3p5UFB1EW8rEbDqs90nbQHwiMR9djRnx/1w+CI/igpebk4P7A9lrVJCbkUl4
CocF5kVSkAXXd+IWC+hx2lRfcB4W1N1x93x7GKh5Jlzdg5rHC4rfqUFEhYQRmmXjDpr6vtl4JFck
pTKZ8GJ3tGpVO4dhPUEMECGa+Hkr/A7/hDxHjHowZLJdn2zA+tDFoxScUAeArzPjqz8hsdqzF02W
fQiGGCvcDptRB5+jKy7JUbS+e5m7n3vGwM1Bnm6SrZM3wKcFiKJaATKZINGSkIj2abAhaGF3ftGG
TdkSeOnaY9MzeBqQhwJH9uaVfq58WcxLZS27KrG3Zk1p+GRD1EDlEpesfXfnkUUlKpi3BYo0eQV3
OpP5IoRwU4hU57M4Jhx8HQQkd9Ng3/UA+V3WkpkLmpoQDV+vVnMD31DDxYJBsSqV6MOVw7YOI6LQ
jwySWvRC6Id4J9FUbkR2CkiST33boTxKu4vjIuit7gj+aIw5X7IePwh2lfNgLiKS6sBu9uj5wrpO
0NDsHq+lyBH149lWwTHDR6XhoscXJhzCjxBI+ykLgyrQxdqoD4Sd/qXRXMTHWIZxRSqxQbc9RvZL
lqH3K31Qys1A0iW3GM2HtIioZImB1WBv933E07mM+F61X0SZOZ341agkdWWv10Ysge4IrvlmBpCo
CTwD8JJ6QqxYso/JtMaPegt67fm9pt8ba12wZc3kLeW/PnRHu/8GCVP0BKxOu8nDKL8vIwoxs75o
M+axlFsjKSu+Xdyd9Fz4tQdlrRX5PoLWt7WdfQICfJHTB/TFySsLNhmZXYOw6BYh8R3lsV2M/wKl
b4ixGqx1canB0Y0SDczvBYlvg002nUdVny0tcFLRxiieBwy8WDpVBttv0Pf30Of5S/nP36JnYqiA
YW7RgynfSKYxanJ4GoWFuqz55fncxHhkMU57IUGIpTK6D1Xt1iTvOx3KazDRQtTB0qFgYcV+dLl6
zg4x87Ekjfr+rWufVp8BUkBnl+4dtfku5UGtvipKhiQnIKobvUKUvrcH2WAt4nCk3JZMc2VJ8+bX
9pv2py1HMPSNhnxQ5QYXyQ004is1HskOIU1YHg3b0p55NH0JQU4fNV3859YY7YgBSx+wzZTdHpN1
DU9KxVxfC/vOoS6Q7MietoYAUh+RZEF8Ag28Oh1UaUNmC4dy7S7IYdSila2uSjsSOenjnXWANvo8
BT6wFZNehyezok6743HCbqmoQ/lkSra5PlqhaMfnYWklz3t+jEV9dCHmETVgN+Q67f9gVNP+xKyt
4Fgm411JSHkdva6g5sjNSwLFnwT0Srcbj+TZlSA8hH8ica8g+awrcJ8jF6dsuF3YqWExZHWiI7UG
8XiDQiq3aeD0GHt1oAAtFG33TfDAxkDc4KUUi2HP559d3CdU2/vTVwBJvnLX5sL9u7gQP4XntiMo
0vjHuUA7o59uuOMgE8FB/TdSGgKQqDro56oz97IGmAVvRb89OUw4gzfcs0xCvk7s6kD6LdE8vaSc
WQK1/7h2Wi+LHGykB/bni5vnLd0b1j/tpMsfp756fW2SRLK0lOCMatnYA1TMFB+Si5BHc9dCRpFg
vJ2M1yesAfxNNuNBS72Yi17k2XuMO1s3RZW+gCR3iYMyZC70V6AnaXuoRl8ZuD6jz26njLCdYMob
ComNUjKaTPmfxENxEohfKqha60sZUCiWJrcXKZxbVk8vQR2bd5RZjZBHNMT1c8sbXosBADyMqtlC
yrsgcINSBQg/iy1ofhAk32QSBqLG3diyAzQ7JdSDiwGKuqAQZpRoxnFCRKCY3fnlL0T77P1TRuqF
o7o8EVNizCxpPDHIr4NDt2DZyJPbzC13NSSQeqmDQ0jWjt7NcHw88Sf6w/k3brVDqqHX4rnWLb+1
HcyZ+iWFiVuqB+buq/c+s6xkHj0JSH4CA3nvHTL9mViAqCDaxosqaZP5vqrWB90UMV5OXiQCDGd3
V8H5UrPhAtJmZpzPZdVoc2KVD9N5K5XY0s1zlFE448v2Lsb/6S5Yn9hj76vImlvp9VZHSQCwSLb3
gb6b+VeufLvCl31z985D90IS+xwLK1kpsPZvmKqQFpy4SLal8+m2znJ5Dm/Bk6f8V2bVjh2j1XRx
Eh6shwnz0V1sifAvVYTaPcTxwL+2UtV1Nu9aS/rEh0attxeAKWVIEdx8UuJDbLUBOO2F3P7FOqHo
RycqiUBQe9sTjxqvEqmADQSmukN9mJGSh8p+wmws18BsQbJPQ09txOGFKlsSSiyLnw4bhn8tB+qR
6mtxEhupA6K5/8Wd4R3Nx3EmeUTBb/AsP0/5WMbAe9OsEz9GoPcSDDFqipiJ2RluGBmyzBSwLUkA
jnPiojfWhJ4SDNf0ZWFVTGzugXTKffeZBQ==
`protect end_protected
