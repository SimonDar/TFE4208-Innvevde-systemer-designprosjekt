��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j0y�ߞ��'DmP"l�8Ws����3#�P����P�ɻ��v�B�*����ހٗ��l�I�$JE�����X�(�>���'v���)U:���si����mY��������f}���/ p�2P�W���v�R�9d��$h�E�o���kI���c�z%�y��	E<|���Ur��~����M��`(��hP�l��	�t�*�v1�.EQ�4�$��f�g�Mty��B���m߽�]�B��+���C*�b���e2���Ab�d#�$1�I����'����[�KC�K�+�(o`�A�o����!����N��a*�ߤ5�Ō��h�����l�fG k�t+������t Y��Ō�T���E4��Ke�`���4q]4�ɋS�Ի*0ט�Tq�/�a�9 'Pu��y����8���]d}% ��g�^��˟ 5�a,�B��&��.x*�����Eշl�,�R>,�6�o٪�,�� �
�����?����3ݘz��?*ҿ�CX��d4Ϲ���VK����ޡ�-�VF5���N����_�����z�K�����g������ۏ�%kԇѶN��4�>��z���T=$�#"S-��mK ��6��I��V^��[��Ք��}l��"���9���Gz�bM�SD�a�yӸd1��-�X��i�N�al.Do��t�8�O�
(�sI��/���RVYi%yy�L��by�/D� ��y�6�lK��%sأ) �1DFi�?Ƅy�}�~\���&��}�=ѽ���;\#t�)2����M� )�j�6��ҒR�r𹑊�;������e���m�.u5�o�����g�]�q�`
��*`DRlh�
J%�dxVg��F!�SɮV�tŃOH��a��gK�|g7��7E㘜�-���7��#÷���SƄ�=G[��`�Ԧ!��g�s�s���g�WSL�=s��k�����Iw��B�'1瞧�Db���.�=W��D�0������.$�]�kS�o~9,���*6�Q�e��.'�m�ގ�d7X�+R�.H�"c��\�3��"�A`^IVL#Jg��s�{t �C�G+nٱ<��{��UuH"�БW�5�$�� ���.�~�9$7	�]d�;��"^�F�
3�����)����-$�9�C�BY�
2��w�'Wz�+	?K�r��QK:}XXb�y�$n��W�V��v��F'Z}�3��~�:���&>ʲ��s����܇B�S��3b�'��3�=^kxXM��B��O�pf�!��G{�t�hr�i5�ش�(����{��F���l���%�7��
f�d��w����)F��i��H��2��a/�%�Vֳ�ҷ�յ٠d:�T)rYN�Rb��Hn^�Zd^d��U�}���\%�,����'9	�?H���<�5��_��ç��ް���V��}4	��"���~J�,���ż����c�u�]����Z����]�3��W�Jt�.�g@�,��;Ys]��	s����!��r��֣F�c��t/���O2�1�c+I34�E�teoߵ�na���{�η������/��΂���&KH�}<�f�́>ʜ
2���H'���h��|�x�3m�e.  ��)mx��!Hf[%�1��V�&9�?S��g�wCֳ>�a�,��\�������W�6���G���M���sЂZp2��Ri��Ɓf�{����3ڇ� ��S!�}�b�{�}C�_�J�������r�B�ي7�2�ӹ��hcRiYw�x��AБR��R얽�a�7 ����W�����a���E�$ŧ���G���ZQ9#v.�#���ٍ��Mf���Ws��r��O�������;��'jFF���UD��v��<��OY�g����&�]�E���>��Lԃ���c��;����vP߈O�>�|?��~h�L�s�z�� ݾ���q6*�:��=t�Tn�E��嵲�i��X�f�]�^�SL�kUT�2~f���/Lj5\�sZ�<���K�d�v{!�g^*CbBA|�=E@R�2����7{�!l֚޼��][2�sJ���]��9�%��$���S���*%��`M�ҫ@{B���o�-5�3���{3n��ރ�|���^Yg%%��>G)͋���AB�=P����.����MŽ���%��ǉk�8�P��2����L�0d����e:Qm
���Q�!�Q�8�T�nƿ�H����É�4 B �*����Ӻ���'\�l�:Yٔ��/]�i�/�#���فy��j3}L�2u�L>a���ȉ��g/���V���M����p@��+��}��H�<��1�K\��M���
��e�2>�s+[�I�r�?��?���[u��׍?����tAu��O臋789�c��>���{}ar�
\*��`l�Z7�Xo�iOs�-ꑲf�%k�ڋ�I\�zsͰ��SH�oP��QTV�GΘ��Dք�D�f�5�Z+r�v��e~MVq�&BQ)��\�L�