-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CSQ05/blkdTocwVPuFo1Xj4yWwqel74dCezy2daGA5tFHoCwQQt42p/yO50ELWU6q0i9ggn8Drg9
rAP9ze+a56LEx8F8sTATYUgtg6gt5SRO9puT/JEDfjeNxS2v3DjYfJAHXYrwHn8T+ddo5sXGv9xQ
FzisHXfChKniCdXn4wMuX2DRfYgzodMvYA+tTOxyCIGeCMnUuihqMEDdnsKt3lP+fj2AVf6WqCtN
Mqul42bO/4cGpKFNF18nkfCfCyCo1aTr+SRDtMvbU3hA3rJvnqsGLkMi4bCK3+lzpPNspcIHi4Vz
np4NBM2ecA12V66zSq6JLbWPlQF8KRZRhfY40w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
3cmTw2rXXTXhXenfYGfZd72fRmYBFKhyjUbQ6JTF/aP/PNUi/EhK9IlTmOWy8j+xUWrEmWMZ651X
CA/S64rB1T1WzZmpfrhEnPE20qOvUkodXwNKIUnioUy74HHWDloiB8T60j1WrlVlsDhfS/ykcPa4
a4pU++gI4S6FoVgXNlD+uTyu+W8bKBVXu/vQQP+N9RH2P4UVe2L86Wuz8GKzCIpFwXznSyF7iQ04
3Bihof4HI49bTd3cQ3ZVyoezclRK+NTnwQFar3zG254lpQXYcxMzjldGKmX4mLdyXZ47ZrLAbazo
SIp2jLMAMFtzMFQINIxL/4eMBzfVYjbuj3jh3dlEf7m/amm/g1smM/y1F+zTL73Uaoz5KPn4cgb2
uJj3cPyBu8ak4Y7q8Dy8rX1FVe/UwjzLl0EkKLqjko6ZEQmNa7T11+juP/SdBXyAyfb9jUAUh3hd
i/izuNmL9597SKGXwMkj8CBQ2zSBvEAYPo2ijWioFWAyxunL/MFg/16+V7whsgT78W0SIDIBX7L2
2HmTYBa/E9+6Wn8/syPQe7JQm48iVzpByFcypBG4Q2AvhCw1iV/Wl58lDq5Ybq6QBoTU38nggxns
c6Q3qgtbG4HC3qu/EnDNd2tRC4J9pmGMou00Wq6t8JHlCkY7fr9x1HOYHCvddBMEhv1TXj5LlVBK
pElzn+TY+ACTnDCs3AYLOe+QdR0XlA4OHQCHjKhHx3p8JgXnc2z5H4mTHQbBIckogn+yQeQsQH+p
hJfNPlaI3KNfYfuws78M7V6YVcMcbV+fKngLYOqMp2qbQOxIzgaNlaFjMSy5qUSwqeJ9hzaHRqTY
4zM0iABW7pVOG6g/iazugNlgdv9TMmgSejQ8CrIO+T07fS+KdMmkSFsbqixVMgs7RkE+e+QEvCli
8qc7XDMSPE0CIkXt14VzvePkaHUteZ7Fa5STb4lbVbESEGQBxMyhhGu3kdXj7NToJzKQ+MmGuJdp
CmNvtPoZ0BWO/Gw0u/hsrWKJOVan49QKVM/PW5xl9ptzTud5zz1jSl0tzdBVHRO8UveX7wtFhM4W
SUKPM2s7KBwJS+UKWlWESF+ecS4unbU+U2X3EkHXiWHQ1fCFPLxZYoHow4fqR6KNKEge3FKiRXY/
bVD1Wg1Xs/D5UKmmRUQYGsGlQztKLccJfBvafpXqOTgOrD26GVDWArlAFTIzGXs0IB0alTVbYA7f
vyW/AlkGGMVKb+mwScVj+YUEGk455jkJVusqjptm8EtqX5QvrAVmByYARaoRqG/thre5ZQmOlz6X
zs6zFKVS4BDlrCBEVNv0B0aQDVK9UdNGCEQwRyAch/eVUJl8IxRqC69/23QVJXXRR0hlx6vMe0sU
RH7onyTP4Z0TX2uRzfdTpqXDJAUxYBod4foJs/5qGce20b8d8w1TtcHsfcGus6izzVA7NEPOsUCw
GncJxhZLzRE1yPJSLTpFPxjdSplc8i1epRMdpSFN0hPnr2Ddu1C6np0gMEyV/bRcto9l4Z+aasSB
buBIKD8rPyEQL7YcQUUxrI8fNljccifNmhlvG0WUrp3q4W5nQ+BrvfAB95999aru4jSOYL96O0HH
SgUfw4Qg9/Ok7AKWB6n6txau9EmdXh/nmAc6EC1aNz42bag2/DwJ9t8gtkZ+glmTZV2ZOrnbavVR
5sMb2s4vgaIT02UwB+3RWKdhyVCK79ALGAX/mBkxzDrMq6B0cKNCo8rKJSDCFq3Cy58ie0bTp5eM
wLj/qcUNCB/xh17E8oS7SHpNPwq2ev+wDQGYLf6GNRCWpJr3wUEHKL9YCjTEP0FWEOJQeVVIOqcs
YND6KBdPuIn+J1Ag2ELKUrQ9KqnRQB1jhSaPHvbuyX4IUO5WvokBi24epUiRWDJqXMxfF2fexA3J
4xPNNBrQnYLqtrIQ39SoP/2k7qJ5Lug4mRnw8ci6vBSiAJnAut0eFxF2yOKDAd6Yhly+AdlBwwtz
ruRDHqiPckp04AkOlD+jwJttB+1sLeWkvnBhoGnBR09vsNeWJMO6csU9gDbPX854g9LwcULb8iLY
wIeSokqEPD6qKMjeHEAVCOP+7hKfquu+sYr50n7zbTQjzuDTJVKhYSvAxrM2rU8P412iO+DzHlvg
/dcMaVRby9HKLGcDBVzoMpk7tihHqTQTfl/ccR1V7NobIhbli9SFY+MX4tXFSF1S9AEWGY6u7cvt
9gsK8+8kOwoxtejfMJ0hR0ZFXB77xkCFk+x1Wj18uEOMsHHSS56AT40R4q0F4PfGS26b+PdDOc/a
C2bUTU9uZf0eRG2uPMCZV4RmOGoVsci1IcIcUOHoqxW5ja/e8yHbRWCnWzhMPGcSOSdzLYC7Cevj
O8mq/wVdQmH4lM7GbtK4mOTuEZsb3osXKAoL9WYthg/rUxJZw91YyFL2sT/BinSvK4/NBcMxJjcA
BaureBmSGIeo3oYHA3/mYmJcMzDzH4g8bUrx0Fs3Yz2ia78jiYuODXF+83SOnJQA3B3Z7TO2578N
U9tcVJ8HRLQv5y8In63aQxm6j+mesywkVAaxFGFGnacoefIUCP8UyB/mX7Ei2qdD0sewZLDMu0QI
OFgHzNUvauvQaX7tVwVznvmVaMLbRqmk250q2zh6H6F29xF00sdE7dq++fLedBqkOVwH2yeJcHbs
MYmMJD94HYo9iON5a9nrmSwzrvjzJxsEP77RJ0C6melK8eS8+6ZcTo9uiGUVgnn3czcAad7sS2Ze
whf/LtKBRghJMJHUSveqXzARB4+IgShfB2bFLZbDgDNgD6Y95FOrSh++rKVSUOGSAEBNTpW4p+tF
2e3U0bz6SB62oiyurhKVm01FPpA9sCyCCGFlqNeYBYACCv3+t7sF26L8o6EW/JZhC6c1QkFYhtYl
0JtWBWsAKSV34IYeV6utZAEp7ny9pCqCrXZli/DVkLvIT5nXQATfQARkVoNyWahdEajMdZ+Mkes6
hbjSD786ti1ZL0NJL89B92feuQ7mp05HIH4v0h4esfZ6kRTR+0uTrT8mk3wKYqwxo8mWFX3n97kk
0rHad7+TDQKbH7z0S+ePXzUeBM8BFKl9Urowvu5ff1on0N6pslqWAHFVlRSSkyTd1z0itIyo86ae
IWB5Zb/KGhrqgfoYqKRIrnc6vUpXDU3xA2lT+Oz5hLkVfjl8PuKM/cOBT69np7nemMX8aeozL6rp
mic0dOW8gcoTquhsEZhR7/1j0NK0W/k97RfrmomTSCMTiouBodmA5XeHQSEDxdIH/VGtn3YbS2xT
dCN4gw/AGrW028y8f8T+E60Cih5yGFvClikW3kIjYgdoxyxEuFBC9gEqc24oEts9koZfTRi7C72d
CFZStl3BSaYuzd2KDDoKNeklhVywZthdi47gFqmHi1qHtUR2voXWhQ6jcxoxhGNBGGb/YkT6x5f5
rJst1Qvo/XsRbYErOTzXpGyEDoNf+yidLXEMkEmgAeiUVhGa2ooaT31nGl/kGAkZAEwwCwA5pDep
Qu/TPTlhzwxuE51R4kUhNSA7xKNqBS1uQilHhoESZnQUiEpRWTnHHCams5ScEm15J0rTGewxAP1H
8PnngwXlt8qNx1mEij3vmdh+lyklovmtZqM0m0PcMjqbF9TKdCNqXB6/r47lVYcul1VKeuWgbh3U
IPdvTKeGJpdyTYwwb/KyU9CRpXDOSW1n4sSi6jZtOcKI16kOvcsJ48d91x1qr/5UiIkbrz9SZrRt
gSosJTWSQgP3Dlz+fLwsencrBN5iQjKeMMaSH61u65P90NsL6Oq+VYXqvxbDgKTy6syyY/r+V5tc
tNCNXRIeRM/Zq5HQ3BRwsvO+tsA73vn8K4AGlTTGQQZAy72HF7X9dA55h27Y12zNs+/tVIHpB4X5
NSOtvPfnNtelF19nqt92Wlu8pB/DuuygZqKpd+I6JADtkpiqAO9p5+wg11EGGVJZwPeCEwApzSx3
55yA2A856c2cINJIp+KekqyvYrAgoBRTtwZ+FA9+CPugSBxhPui8V74C0oFR06zaAOLgM1aBCau4
P873ih1WGOdKS3fu7ATCktvEQ//D4YlGdaPfZJrS0JgCZ15m6Xh+OUFHcgalL2Vz/Lo3P1NZvNqk
VMvaBJ/8WqvZOqf77PcP4VEXDySMnKe5LDJvSKJ6rTVaq2umxSUtcJ5bKhwBX1hRuqvjGp1wW3US
mPRAaeEeJWA8ntTJzI7kZmVzVd2l88POqguSPbLS974pgtpaYsXW8SlMFdsB5p08TjKLx4lMPCJk
Z6gDy9pB/BSu5nOGafVycQdovYk6qq0mKFAptQmsjA0z8wnqs31y4akTWZQ4Xvo9DhmSEIDVSA5F
cZAHVrMYpkydKeFm5LWeEIIBatwUTghUjWK3Q7PoeyD3jZJr3zxSsFvjwpwC/9t7wQJKMhRoVzVp
MnZZH+whr6PuwVVf6hR7KAFXsZhIA5BEC0UUhWwyYQp1XpuYJHcAE+XJydX1RxoSpya9DLF9KPEP
Qikj8euQCg0fGOe8EgHfOnwtgStxpRfG8MO1pvHp9jtROPArQFpjmalxOZPmCa0/7U4akkbHHfGS
gkM4Qj81RNxeHZ91VABkMkSy+sHOyTO8UHT78pARY9lqCnvivIU+udsKN/f6cbS9TxOu4YFxw+Zv
zl9MrmYDEgEQm8t8J5MCCtY4K6/gnkqWnsGSIWsqSPu6k3O4vqLL1vZdUoRFA7xK683cR56wLwcM
8/BE5pvVBOsX+R7jm0cP/7OrOj76IbwoTUbHYdsYRfZNNkR+OmLX+sVTjNyUGvKXlHX/+thQRIJ2
QKff/wg3uvodWO2x8MVSwWbPz4RBZsVLlG9Fzv/IVD8P6Vo+GpHBkGR+DJpB4NV+A5HyJZpaonez
BnJCCQqAIW+DF6mMbxOVo++QH/YvX8JyZuCfdsnQssgpu6SthG+MXfpLEcSyP0MYePtTbHvHzzTR
roTB/s85RYZYCHmjeySAmO58MSCEXpptouDL4X9PGYWlmWBZB+13rh2dYRZLnX1D+MI7mfbAYHzd
Y8Ysfl1Tbx2cVScdOXTxfRVePjutuAUGnNe2a1yMUXUufxNaHZ2Fn4LAwuIAC6diTBoMescvul6f
p9plUjyouHMABiPCRRVkXDbajWmLqyXGfGmzE3o+BkxksYrdCzZJbKskjcDR0dju5jkBLxD1rDFD
LetfSEx6lDXXHr4ZY24QylZyyntrNU45zHhsTr8DqKXjsj/y22q3IKVCLt9Ck4mArayo7GtFS1Hg
Iwa47c0Aug3EUlF0JgWwjPG0FoIwyZpltuphInUJjA2qMAuc1+vk73INP8PO5aySC4OEOnq/s7HJ
81bWOd+vzZZOoGWXuGl6Yavc3LgAeprW85xKQSFqoBSiXUnH3lcIl4ZXdMJzOjzo8kQ4AvF9+dj/
UFPE/wyuVePbdq5W9qUIc8aVJTsnThg8YphWlCHPf2+8mwbCKxO0uAqnCa43nRjCtWGd7BznUIu/
fBmyt+EdviA86QFtWWwfwt5/Db0Zpn7Qo0h8Xg1UBJieM2iIQgZtvexAq4jsu73iU8hCdQ2uG+yC
uQU2hDogDj0hZxuigeKzow9kMFLUblNkj1OIYqYNuPXdFwCtoxPy9x8IoUszFwda9rU52UF2GquK
/SSfCF2uJL9O+ub1NK0cgX61HKutC1odM2/Kmk7X+2xqLbQ81LXmr+xgM0uTzcjZKwU6vFgOk/GX
Og+i7hazxZgQMu1RtGLGq/T0We76CSllSC8EnPFTfTiSvbQh2DyjNexmZTEYVOMQpx/ZIHqURQXK
TzkvO3bhZ2ize6ICsAW5qJzActgITVYjS6SNsJ2lf1Cb7eitOAN9FlSnn1eVyMoNoFT9gdzujcV6
HYzBj6PB/ki9YeeCEiYDpMesGQzFCtgEsZ1a6Ufpq4EzMOFqCaaGDdKPe8IXUIOmwz9HGrj90rzd
phEdMBxo2H2lbR1ecsKRjoSlY8a93oeKQDXWswsoNHlU2pIlL2/7UNXW3sS5FjkUuTS/eskxwlO0
ZW+mlBU1DOVfyc2yWDGGiFCy4selXJjcjfVMlOnABPmaxHt8EJxHGoRp04H7oCTc+6HlC+pokTYV
iNsns6TN2YsO4s7oWuUbWeliy178WdJzK70WDbDpE2wHsfVZBE//VmpwpnqAmQ+bDtZKZiL7lHuD
PjMIjKTZTyoALHWeVZMbp/yjMUkKGIrX14fYreB+KcTbHSH0/+vjjurRX+GM8X2dUTHl6i+dkKbU
sPuqVqT+3V3bN03Y9T5ETT6MX2De0sXCM8/wUS5x7DoSIeOl2U2qf18QrRau6wAShIEZ8fF/VooA
1VYhhjtZSNQpHsnc0889cvzKLVuoE9FR2uen6AZEVrNNYHqdVUnRfueEKAFsXLgw1B/aelSPcLuq
3m9NsUY61hlIfwGLTBV5Swm2HS5ryRVmwskx4QDlufYCAjqoBgeiIzCzBTk7A99vSDrwUJ2An2NT
d2wtH06Zt+R0xgc5wm/TiSgv6kaeaWbM9/385S937QK9wdy+gEZPEUq/kt56N+H6ImnHFc/YOJET
/FFuOC+BO3c7HVuTNRgkXgWzemtR75irdXQGCihLa7tGM1vz541I1wtOA6p1DF0N9z+xQsbstJnw
7E5q001cRmMJBSvZEdIuvAPcCcFnivmC3mqvk6qB77uMKHIWaxs9vTf2/IBNz1wotESlGyCU2nhi
s6g2db8E267+zKacGyiDrapV3Qj2uAcdCy9xR5IZ6rffqqZydVN8/sd/m2+auGzwblDkuNgcM7/n
ERUBMhO/tH0rGyXyJBThFYsQfpEsG8UI3eeF4D8x2giwQHqWAAGM8wdTw4m4s8CTexL6e9p3VfA6
lzIhHxWZa8RNR45sArINMzfuE3liFlzliF49hYoPzDjwyhjPHXK3XogusKVMBaeeCi96UntWCAjE
8D26/hGJEYxItZPOVz/zIc/XBI7Y9DBxNjlwxsEnde5x64nf5DC3XxnLuoRzoe0nFAFxTvEn0YJf
IVB6b8Eby+L2PmHvJpvBSWiPyoEhrUEvka7yUPjoq061PY+Sr3lS36fTeEbk2lp3l+3q14xXGEwj
eVPFbodr+lJmbJb5VjA/wWbPgrh04sV5AjzN9DWNH/I+nKL2oYUwUZEFlxLPD2cefPMhkG5Vgqkm
+IFD8rEh8FPiNWY8HE4/buVp1r3WZ1Qu+fd7qws8LVZFVVcycXTACqWGQ0/zNocSQJzUxflqtlsm
kBXbpEOaUG4cSu60SVX9gm3TyxLym4bHFhOmySNcQ3YLqI82ChMVX6O5yB9BRihXdi4loRwEkw58
TrUIFiMMKepIgsce2kaeM8hW43y7WRebAI/J7HfoMaYPYAE2G4L5NCpZGyptUaZPlayhr0+8VD96
sW6W8Xamwm4AG7VJ+zHc++NmekPTPWyKeXVaGp++nP0VyE1+tq0cyq7aiDbBf5Ud10a4lAE9TgDO
RPdB2gdyuzjpmiTbMc7v0a5BaTGItWiKdqe/1oJAaS3DGaPoFIUMR8tid7r+IS8hVbMBkyJIVazv
ydjtH0CrxuWx0hT+5tMAqJm71Fn2XbHxdEBt5XoTdkCTB2CLp9SvL+Z+5wniNKLXnwlsJTxbFrPs
LT9+NPKwopZu7FiMDYpJLmZYBY+h9omHy4+J6VfGBPyC4z+8o/FaQouBfpWh+who8ir0MH/nyH9u
Cv99cBKDsMwePIrP4gg42uPIWZHquH7t6yDlbZALkVZrk3eY3sHueGMkPT3umuEYaceRUMrQCWce
dv/E1q6TutSr+s6BDUFc2iaIeNtSzXc8McxI/NlAh5huu+q/tEBoEYuF1eGiBUnIT9/d8Qg4Rk/b
Kzw5xNMAnA21ym2UPeh+4uZw0yvw/gRG8wfweiMG0BLDswUcktaq59rtiQeLsHiaoYNJig/IXd6F
H4C6a97v7uFyfXJgl1bU8WEL6z4KyzjN6KIT+nr3THLiqNvYXcw1PGvoWmLlkh/UjOTsPgw3Uwyw
thT2y7kKbh5JFYJkoRRJsX8S9dDqLEf9XuqKuCQ4x2ZkF2W17eb9iG0kdvAnuzwGNp/0nR0Rf79u
Emo1tBPQl6RBjaw8loy7Qfvc7QdaCTbnxqI1Yqp4kO3vjNnb/ZxAVAPpUZTp8FVkWGwyz395JVgY
j5xrIp3r8HkoF66AIb2Xw48aVHjUuS2AyBgPEecdOkCIau1kTtAZPFjYoygeHsEdg+WXej3AwPnU
iK0S7Yx7vl2pMYqvURpW7YTWtRL+kBjb4OYWwCc90I9kGzrXOggT9OHQ4EIoz6Fo2kZ588YmvIBb
y/3cOM2g2eiUMEX9CrTiAulc2F48cnNetu9Is1UYKLL0g8WOkF8rCTrg+DCc0KpjdQL4wM4SxqEH
aw/fJChfgrFvAN/oCtl0IcGg9T7OEFQCXHlyM2kT5QSIaMdYiU2sVJ3Qc9e+HOCcq44SDg1AJxYD
ojKxkyE2UhjmjYWnXZE2/VgciT1GsoJPFzw0eSHfKiFXBcRJaGbywakKuPWGjJW6FK+l6aqgEbeh
pfPPqrLh5j4JWcH1+2L6TTQNZKJqVDAyQFFLYqs2HFiMsXElQzINJfgniqUlRobe083oeR1cOU1c
8PTvVGT98G+fr2uewev7usbY+mRvJJNS08RRUpqaBMFwqkP9Xjwe69XUjDQJixkpCcmfmeDlb5U1
GxPAc5ERqH3ycPMISZcoM4CS4eJWTSxbqpVulSKnxm1tG1oXpG43XUk7Cij9a01kPbtZKxwBDBoM
kbMJ/slaPzrPy/lncOpbQIiXE32ViDNz0KjpnuyTEDYAehMgwWiXergMUNHH2R/9aVRYhKAoGmK9
zVoIlClPWiwFtgDJLLLPCcySS0lgZaeFFe/PDrJW2fiktiKla9iP7/3xRztZHyk4ErHqb+Ea7Is4
h571/B4V/JgDsWJSI8MOhxJlL4t5AJX9NED/UXJhlxZk+X2vALrjsfx4bJB/0Ol5Rx/dqNl2/8N1
r78ZPYoaFr4jmuNWksPVbTR+b1pGrRXw/mvbXHGQ4Xwv8AvMbrigQVHhLoS9WITlsKUguyQwZ1IU
S7LCAutlT+tuGp7JEqn8u6ZWBewVU07f4P+jVb2BQpvTcybUKlHIpGA34gHGNz5AgdtnpdFx+pvM
n/c+oFbOfKVws+pf1gt+aYtSig6RM/YDGhku2g23fd+UIpWNKaos6fatMH9ISnQwZsz8pnqn/3PA
5Gi2hirODK9prnjgHjl/WB9VZVwaIipKwepBJL+uok2/shj7adSGKmmRq3yfcJheK6IkN3xJjh36
ODip3bj+XI3dcMf2ug4NwFiUWe8x9qNrtgpx7w95rRkJVZTVyKwgtAJZFADPl99cjG+3jN2BN9xV
VMANZ7xMrcXAQYp3DXb0KsoY5+JMkXvzH1jsevtvqduJ93PAZOTaQgZkRJiKyAKyl9VJQl3/YP9f
Xxk6H7dOhRsrYyrudab+QQODje3OGfNM/NHdjN6/y0vOGhXsvDsVB7VlbjdP4iWPfWmRmGXl04SP
iN7JDleP9joAPvVh40oXFua1QI7D4tjE8eVZfd22lw5XWiy1AY/3ZKzB4ns0wtIXgySn8aacOgjh
I/uDG8aaEF+oUn0JBON4z3n8WDBgEXRzkXfSsxjhE5cypCafwHU5DVCVgfDTBnGVFjG8+Uw6rYnA
9UpoBdLZycLhm55lAXat29qAKVIm6h3kO/f29qytyXU+3lmqM/f+K5OU7IQt0l+03f0pxziKqmhI
J/BZAQ8f713ZNr/jgP0M+5MvWKijTT4QKZBz9qiz9UW0HzAWvV52q9AULYRl01wVXQ8a5Ec5Oeda
r/I83kyz8ilyib6Sl6sBEvbG0UofQClnVpPkVZCs1DdUCz56sRa+sX/xDHtHLcsDTqolWyKyaxp2
9B0zOETMnqpWVbJGIeC/J+XkhojGQlvROjIEa4zy7BwRIt1wR6ac1ZN7NpVmX7mYj5ADL0yEju8y
a7bMLhPOmweqpsdr213fF0BUh79AMxZF240eBQSfud/ZlWtUX7OHUAmhYZ1wn6IJibVEDSYkekwj
Fa4wLBoQkeDDhycHYliYyuvk0AJzEz6AOOVmnSyHzBwHOCZnotRPYQy2faRRSLFIcsluSQsewHac
4E8O9FIetBcW3inx9sQ4NhfOOtdvZFBt6FWRXyfVHa+lyoT780uYvhL1LVNIH22aRBpUnzr3WtLa
aM0/QaNv/e3H8d7G781AyFyXQpNphRbT+zFAk1pU55xtpfgfLZYOuK+K/jLZ6nN2BwDAbCXqDUzX
wY9rUCuiV3CcUieM0ghckfD1vJlYZhFDXuUHI8AGXYNby+6kNboY4Vb9M5oWbZAJVLt3UwAWFVFu
WruCHbAOTMO/gQlbQVKhea7JfSGFqI1iczA5bqfWgYEgPS8pfY9q6T3+k3bwyqoum+LWVXXrgmV5
5qDB2G1eGQuzxowdOePHobQskaB6L+FG7JIMJ2WwRzsDxiyHRipTThhODr4z7guUukLfrRQyYqLJ
5YrIPY+pXpwiVUOKREUGKarDs8qDu+baERC3ZgYuWMpWf1uK4n4zqwxH1rvIjqgd+bxNpxDCrKhI
JpqA5lefdN24SyMK4VYQ/EtZJynBV0ZRB9sVvtx4aXo08mCKMHIzKXhaFFv6sSOavdMSEq3sB0u/
lonj8DQjRcsKVtkckmqKfEvPfPo8eHgkqqH7YUy1+T1gy+cFLr3Os1Bn6RVssr3Ky3SN7qYiIiA4
icZOXvNwcZSEUtCdnHb/MlbzzoUa8VAaCmVXAz1sdTDCItY0q7qvA2hdYkd2Q/l+hYbTQeh5otum
9AK3or4V/kISnXNE4bfeijo5dASlDGRwqr6uDs7LBsDSr4SHSZudDfLiXXu8SlhT27Ej+QFUSyJk
jtamBiD8i9rVdYkrTdbUyYuG2pERkV6C/KWDp8jpar13CiyvYDBF41bbEHyLFNYZiHuyGzkfaFjj
`protect end_protected
