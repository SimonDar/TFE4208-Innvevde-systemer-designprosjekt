-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hs6YXRl6bYzYlyD9gaKmnEMTMBIZORs2S6WdGw2VJkHzZZ0wKIL12VX86TREd0EmNsyaN72TvvjM
KM6Hy0kW3dlhtttDpTLqAtyUMalCPlOTs3hIq/ZJzriy6PC7/PCHUqmj9C9m72Pbs17EnRWi68LX
dfC85cQAEEo/pUASpZJM7AdWG7uHYG1m4GPlLdCwtkhg8DKGk1NE7D1mX6fFmemaTklkiTtC27jG
rznn2NqYcw3v2hPRFItZ/qCU+a4cl35UavA+ObeXsGJ5dcqEHul7RF3ghQmTqd+7XAopjXZ0mAld
G+hde4kZK34kjQG21y/929CJ5DibG6kySQO2xw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
meg75oKz9hrGgbLRvy3aY9PtfYTDBkwW/n69X6sasCRSzv9Sx3cXNR547gcJYgyrIGnn7ZFhbynV
eaP0ZtW29/KERMclleyFoDr7No2FJXXCbHivG1GqcGlQ+47434QCq8VA7ysAr8A5gkIfEMwdK+c+
D/ed6ByQtvkhhFAPZZbsvmhjvTxIRK0BV4iVdjO77NikFu+B89rP9FbHSEcJMmJYRwa4V5XM6BFS
OuozG3jjTjrBCf7YT/Wuuy/di+yVYwiFBU3LDQ6HOe3QnApxAfehjzCztzfYbuDeiQoROHFzlYnL
PjhvMSInd+oxo0JzQGREHohH6x2m0/uND5q2qXjH5PkTkcUGX/FzWNhHMenWohtWWQbSpZ8MSZ6A
rJkgse/izx91lnq/YXp93Be/k82nNg0ktKUFabOkNlxujiaC2VpbJOFkQzuFoDL7ZyVBRDXlBHXB
c7jvCF3VTaftLJLnDrR/PDYqSn+hnPv9bf3egpAdXfTFpaoJruuYj0witjJpmmMIuCHKAWpk+JL6
9T5LLW70uXPw/jm4yfwQpiIJP6asbpUIYzs7+mPky6Th3H5gdGU4LyRohA1NjFySDzUD/FVp1/0i
LKoKQHsUuJo1rPa3BItfzjILS3aj/rUfVsEQLV+C1N+rIJ2DaKpvDVc6DCbzeECp4t5/9cNSYAI6
NhR9tFkGnvF9tRbXzuRX93hC055CXtkfsIxOfzXfYQa60kMNtKQV7INZb3BrROJpwRZ/mjKlt37O
cU3Xhy8aslKHys9xdTG4AJjsboZ9hjQwsoVBCJNfIFxiVf7wKn+i2+HFx8MDTLct0g4qs+wlaeZK
7tH2JKrV8eHJcmKMmuhfLtGwkFdcGnAFJfp/jP1xvv9yH1zihYEvnaukRGc5zxIwmvVnSxOGncGV
nR2eODxfJAZdozkLpwx2PoEpvZcIST9SA6mrJrMR9zeAmulaq9lwZs8IFWbQ0zvFmtHZMVmHqNSM
w+SnLbl5AyTvoNcbCBfN+uvDXYcK40aEhSJrxSv9YWKWP3FryrunylD5nWMLX8BHK5b+eOxs+EqC
iTEG82qQSVIwH6hvAmdJtRFqcnTiEzX1R/WqSCxrjP6i5izjhqt0XY2r8Ja8fIfl62uQEqPCmEsn
wVWdGTbb/KudXM9G3UuomKAUH2P3ARthW0yfWbFpbuui0LAPKF/iwrCW4Etztxedn4EE5VNfdusX
8HM4xevIhkbcAW/Zh+ClXVRU8xEspGI6AbWiSIGbbHl1gbJUIzwHXiJfuLtsY65eq8Of/XmZI2jp
YqHsbkSyR89VOBjoCnA5X3Us6l37KZmswIf9aDUwITDt+P1D3JH1MRZ20ni6C86jAGC8qrVFu39M
wyAquqQ6goZ6yFpd9I5uCWDg1Q0wu0gfLgO1+9t4gleUq9sv8FKCGw0+BRNHnMx6ntTsm1Fnk26f
4hTpo1Jle2uh0iibWlhjW4Fcl+eEKO6XZY6PQnPvpjHGyoThTRGvunEPClOmIcWIUtXxa9C4MYGs
YzhuOh+UESeMimNReto6xGFXfMnQYqO5ZgBZVH7fBCpCRUTZzSdQ4onsyT9nqCmsdFo7g6TYbsgt
KOiJNdnFRlbqXxjiFpa6AUj4ZEmUluCnOP1EkUO5B4g2YrBzkXztqumSKtV1cAx3HJ9VJ/VLFkwp
41BY0S7x3GmV9aKr5aD41iNaDDf4YFYHZKM+gQmgawpmSXMe8RFn6wqy9QoNiFlQeA9vYVClE65a
yHRnXmmBqNLpAHg2Ss6EOyQFKKZCZepbzKnqoDhSH2Viunwbn5dA2aTz+KuahhNIsvT1MHFLO3e7
iD/4mO6y4puTXbnslNHfgl4k1s4yQSiB6qMSAlo0+wFJdSpGfr1JEUlOmZVjBxV4Y1wCxy+7sNTJ
tjI1pARXbvUjW6iEd5oRmpAyfAPKH6/hmTOfKJmf6DBmEUyCiYQ9LR2eswH+GB7fNagiL/Lj0ilk
A025R4Jx33+HyCdnsz7p3LwjXzV+zwGnLNRX04yrn+X2p8A0ekaaGZ7NJOXzySXJmtUTp5IEEBQT
NLCBdPEVjvoct0zUtW8yYBI/fd0EKUTKIBZuj3uUp0T15x0uiSLk5C4kY2Pih+4AGhieLpw7wtpm
2KHpr0Vys8h4ohD4N/EDL0/3a69nJhl4oSGGDPVraG/Y2rmZDDyw3uSJzoeBFIUiKTmfMg1g3lWB
sAZa5lAREHRIDfqCcbAo+ZthL+KeGyyIH3PHDGQwOC4PDxmK4EFyAo/7RohOVuf4gsnp+AcyNOVU
EeYxoKdkNQcwJJbw4IpTr2DE8JaczdFEgsRC1wJF19lDZj8bc0fKfIiiusVtpu+yVVLhWJX7bz+K
tlHqfdam2E3C5vXD2jrBbTsm3Ax+1e+Jg9ozTDWjN3ylaQbT3vrR34vgVS1S710ktk8knzsi1+SH
A+4nM8pVQIW+AD1m1MkJdkUh6sX42hCSmkxF81bJmbySp3kY5v3b6zqOCQNJfBzl0gr9g2z1B/dt
0LbmNtehWcygI+pIebjwkVts0GzD5eojjTXYsosa4SCd4BIoDE+qz6JFy4ZlyPTmAmJ2rKHZ0xnL
fjmf1+I7CFBLFMjyrtMvWI3UGEfGunM8Dpxmx+dfe3hWWEO7z63w8zEvwf+MsyKLhMmrdWyFiAcw
bSrZ10JBRqyw08Mqt1H2eNjBivZwIYFQ1LCqKeugy6I5ayX7HE/Ct00uzsSTKpYAR6SCQF1vyGHH
VSivkOTTLLoxGOynX5j66vFBu8Y4XoqcInPBmT8979JloHhKZ+qZCJpn2yPRfiHLCNFOtm24Y+Qq
cqPFvohLc0w3sh7BoyTLcG1zFCbBKVfp/wVlj2D2SwEu86Ge8ZMcEL7Ksh765/ny+HlaDTwamjQu
Tw+ZfBGZsBwEOXVBOzU9v8t7ctoEEgAKTWtea3SR8+f/S1WacbfOOXWnChuCJ+JmnDdZZOxi6AU2
tD5a4RlPWL1PaXTNkjXvtvyXy4dMcwD3qwmMfnbB80H3oRhnMXFm8nA41+z9+FtPa9ROD3IUHCbA
9xqW1e7nlWuqEMmuoyRhZFfPfvuwegkyqqaU9dMZ5yIXcBLfeFzO8U+b+6kDsrkXprPFSY56Usmv
PM8p+pRw2V+5XmlQR1kBiFCqSQCOmeIpYP2aKajvVL97cQuIhTNzUBHC8GrqnqXsQ7loKP5jNxfp
gfX5SvbllErOrLhzoa0iULrjUgbUnAAaBHJB1POXz6ueiHT0kJcwdlsHXFzs23q0XZi2/ozoaQjk
e5E7jmaY9GZVRUROo16X4/VqHLQHwrWBUBBOZZ4jNmqNcgRgmD2niMuole2ZI5Bv8psk7/Apy1x9
l5Yw7afuZUWRzLO8joSJqOHEZt39iVqEe2IoWcZNyHBbkHhRs9G2v7Q9FzV966nPwwBK/+bGnXRt
cPv7qR4irt5QaRy1o5TuxlaYiLlcRwS15Y1DwQuiU0y/E374lQj8lyqDnXYxiwsy2zVvWEC6e7+t
n2hyMYFeTn8EaG4rZ1PAE2uVB9OBrKAuUSoICX37qDDIDQqeLvKYFqEmir1xLmUj/wrha1C8QlUs
09P/LMY1xc7iIHAl43bDPBLOCfZrrjEP98QZY/v0y/QfALMVbTYrsuOaYxVhIHehaLWP1sevvNwE
a6OI++Qp4wlYtDTzCy1pW1IHXowmuOTok/7ytRwWsblV7psX6+q1eE/fmL6d2Uz/K6uyWGq5euM5
nk71e89vY+eTAzIPArunTWOBZ8v2/+X18drh/lwopygiSoD5w7Gb/Hy0QVIe28GsCM4KGoAOO+Ei
GWSPmzleSKSdnDeeXg17PY4c/+jUhs7vkaFNskeAL0dciqSfnPuSclchwFiaq8lCGuBENg13y3Hf
At1xqdYziyLAYaykHSdHNmOgesNkoZQ6KlhnGchOQz82FiQri3ejOx+wsCMSHg0T0Fraw/Pdn01E
fzDT78RFm3lTGjQab5MK2GLI1SID8bKkFhFw8qXpC7rJbQH92qWJkry2eCiA45wSVDOnIcsPIg0/
583U3avUNJSiApIW/m0BXdrD4rmlQsjmbkY+Q1S/kaA3r5Mote8771qBxyh8Xet8sNDIGTBmO111
5CvsdAN7+bH2uW6ALF9phAchKtkAV+FapOxagTnixVY4zFLsjv666qKhEfM7OXYbjX9kOgmb4xPR
yQd1F0COvPGX9Re30gpccOxE14QQEI05CiZgSoGToTuxU9dnN6sI71x+xCN57L1AD7+sAnZHyrye
gsaNgXT6D5GWApjiTJo6Ms9hs4GQLFCAEalU5puO9ksq1eNUP/TL7wo36g+MlS2g88um+S/YHmy7
FDiKK+9NWFP/Rt5kD0BKGmEh7iTykyDUEqf2d3WYFQDKCpQbDR1UxCsIYygZhRB4gaD3G3jtmjWZ
jVmtf1Dx+JiRoQqM20E0TrSqYLGJ5xngO22Kvce7YPsbYThTiZLYpAyIdazrX6oqOVVucmxH04EY
XQCIF/2HdeKW0BVy89qxK3TiVIgQ9AE8Tgsfrfvua5BoorXRBRDdw7qSaON6i6uv3UYmqQ2iEhkU
IXN91GLVQEawRuI4LaE0CAlqCkbIAbwXHPkPyUdC9o9iihcnvc0ZMtyLSvOvRpuOPCg3yYKEIlXY
i04p7rYsmIYU5ylx7qOtKJrxSXdvMUo/X9U1mC8L+JgxVGtCgHKmgXayDOPZx8Cor1eJ8qm58aBd
p0McXey0UYI3gx9HwsDr5KiqoNmNpNSsVCbkyIdCLyRSC9Rp7YjnbK7CHivyVWHEdbMJtNi/G6ZQ
sECJne2T8GaqVRudvbsePSgOdhHFFw+WvDhIB5XTSWQos75bLf3oXTNBn5bbeM1op0FD5UzuYRb+
uP6YOFHXLT2TpGyhMuDomNsMoo8+2i9fabnyIp6I0u/InzQeYgYkYSfbG9Db5cZZgltXf8M9bJne
qqHJdV78yiomZ42r7ExrtTEYbEgqUpFqpQvujbs4mQ0hbFNo54rE8HkWyFYy7+rFBBz67oKWbJEI
RfL27RTiRsyuNq1/JgsIvlEROmoNd+wTz1JgpGm2BPbXYtxTdFd5S2yKCTDfstmcm+GFIlSEhxpX
anyw8EIG10GBkuj4ChyeY9BtCA8qv1rbXjLxjmyDHsUDCcvEx00xd+gAqHGmH9Wj+AGDBSSj7eVH
KRGCzBMp4S+m3qj+fo0l4jeYoprldJmULrJOkKRYxP5FLrnGldih4Fc/jgW1YXVpOY6ouguTAIFS
GJM3aslFxh1Ulle/kEgoSCzqZB1sUc8aYUXJ4pOhVRtZLiasdNd7Wj/OtwEATgYRj/O8SQNuG5r7
BoWp1/MUnNFUCDJ9jhrNGycmNXNkGF7bC0uZVOwy0hoEEq9NA85Zf5sTAiEaD4hRGYqUbpwS85h1
+Kti1QqTfaABEyCqdOqxxVdQtHARAIpKzrlaMBFk/Ewwb4EsClV82CxEmJNYQtuVRO255YgEZfTn
x3XKiNcn8VzQz9KhG1RWpY33wTImrhyxPbQkkDmM4Ikwy3wHDVsUYCGV7L+A9zrJVUxhzKNVZLBC
UruGiKUXpNdvzmYfkIh5zv1EsoHhAbbUJlN1j409dJrPlN0SQSWX3SzWzn/RGJ558jCTbUm+98Y5
t0f94HqLeEt7wgK1+NdCrcZf3kJBQlylkEyazXsBnj7J1I/3coUASTe7v8jmD5SbjowKHXqlj3Wp
EutkBsnpoY88u6hFZ2yLozEf9UFJnX4MeZWbmT/Bzjzu4dyG5xUf2Nof+wPNXQ67H28TQCSNiNjv
K3e0wB5Ye2Yd35lRgql3M608U4N8K2tePnW2fVezae1soshx26gpw2JhkkI5s9iVM12jaKC8TajD
CyEyIbQIYtJqWm8Zt9jMfwJwGRLQaJ4Czv209cOXzcNrsurcmhiARh6O0vv/7vdjtx/rSlVOmlGg
j61easkxm5pxgvPoma+UHfhs7ov1N+9s2pJRupF3EF/aReefj+OKrfZT0C38luyyX1YPu1WpF/wC
ma5st9oFc7dBVXc6Zoy2Liiqrhci1IeXU8gFsb2te9pWIOGIXPdprgJiD9W/f0Mgzgil+7vJshjD
sh2b37EW44i6waTBEHRFegpioz8tu4SW1CDbzqB6yepR3CAr6JPSXWMAaqnCIrwf9vDz0Zp/v4BZ
OTH2BZynhQD2LKbn0QQwh4cAuO96jRlce0/7VCB2g/nywFUJlKCNHUurbficfOlWg/jfVQqfTRq1
zaQo2y1EevOh9nf2lzf2snpuWSFvVVNfZy9cpyceDiMi4b9nCMsWnc8yOQv9Y7747NokiNtrtQVB
jdxr5yznEHJ5Qg6vC9YXlfjX0omEtHE0civmNtS2upAjI7gwt4bMseRZ3rk8zwZks866Aq1UgXXH
ykTwFRh7eLomJVrCuMBSzL60D65iiwuzx7k7fn0YcKcfBb5vnmU3nlfhziL/9Tn6uI2DSkAO9LXc
McQTr/MAqTwcwPw6atLBsf959lfVlhHeO+aeuihsyKROQFR0uLAFMCJc60u+lLp3mWDuPgCpgQ6c
a7PZ8/GzIyiLC+Fk35WPfaKPW0AgE7JwM0pbh6F273QOYw4k2FtID3OAY6aIA3iNarEoiEligy/p
T628kdeJiBse1786LO6P0jZaQWRUf32TSZRbrFasKPi5PdBgPd/AP6E+iurjo7zjLvzSLR1gzNS3
IPQxiL0pbk/HJ5tMJeih6tQVMWRF/kfmcLdKM1CiOvdWCrH17CB0DYlbi6Fx7LKnvG9veg3Tl/yb
vA80ECrXTlxybSi1oWuSjnVVHMcbrQ+4XxEAhWLWslZyKdPoVPfcGEa7Iqp5orpHN50OeRAGHfHO
yZOHsw4GO9X8vlovYUYzhxUDx8/LGqkkm/L6K4JwAEF+HSt4fMiFIBzPMRruVhPbK98BxoaBNWFe
5ayAw3PI3a9uXpJZ2Qv8gpKnKINMCcYNua/V7iKb6mbFC/gjKV8vJB5Ec5KZw4/mIMJHzrGeANS3
DsNGddwJfeXu4hr5YFJJz+5DIVU63R0utTK0ADC5LNRlEnd/3+w/r5sKXSaEzDaEGFpIlJGIEeVP
txBzN4wyVR4Kn34ovnpQmwnxiDhslo92DWj7evyEBIOS3v3BnfBXZz1iOuWrV0VCUgKVhpOkm2w3
UrNJ1lfOgJEKiQ78E9SttNsCAqYJdaeM4/DPsbu+oemID2KcBxfplaCJhdxX9hJk634XO00+aUDl
B7Hx0fW3TLT+jih7jcrcNjEMACQ7WptvqiHckqOD+C7pRqgkMvJSHRIZnCZ7Tkys9DsZVq3zIfkZ
nxF023vc6tYQTe/tEjzOjurvVydmf6KBUdImmKrDG1ie3zRV0esoK8qLlne9q/VZxmCYcsStk7HI
V7BG+1/iuMrHQKRrs6FEyYr0Lkr+YYKGyntd/3h7LhwKbV6eDXHvH+buJauVFPSingDEXHNQ73W1
yReWOmuGKoClJb+lDrEpSeP0HatfbSeRF8XLHGrhP9ArawxCI9wiln6ctOiFe+A5ma1yuqjwk7Vw
Ye6SXHkUfnuhPbxaUslsRaN2xOFxi2BtyaayvZQcjM6q/RiiHIWmU+OfIYR/JWCbC5JEozo4Sdqy
JuKpTZq8FkOT+LsnsfhqP9aoN67bjn5DjVD1LdKW3VwU9bIfYzVNyeNhqdnIQmCOy6obIfM5JWld
+vLVDg6J64agrU0cW1sJre9fYRkpjR1RW7kX7d64ipABmUKirDf34pcwLo4GtBUbd957vl88ZojM
y8wdKfMjRO2DtOCp/69K41LZVrgljBq5Z04m+jmAo0ozCu+xarK2eE5ZxChOLoDuvuYIuCpG3PV7
fD5fdrSZJ9ArVtWr+hJPd6SnoL24xSkUAjYZ0tiXZnQdL/xtezc11/2lfTKrAxVyqAETJuzk1tLI
W2ID/5KrV6ohWlK0RZ0ComAJYVuC2ssbjpMhTXzv302CHsXcyejMzUn8XkupNH6QYKl2lPV/MPz2
1d0ZCvk8RVZa2BgZbuRowuaQ+GhtCWdl/VjdlK8je2q7Tz/lCyTWjuYZIDhgQCw7IqMaFwFvw8Qt
Ou59Zp9t/AkQ65iZn/3YSZ0LxkvQpaSIoZQEmNuigTsuYCfoJsuTNK2cqlflLeLMsDY0PfHeOTjL
oeoD1VEUnEH2O9MU3S7GmYKBSvElgXfvtAKdXnD7Rtnj30h8AiyIizVKSp4+inSNRklPSqXAFNeD
9k4SV9nw8rgKDovgPejP3OlyaMxPoKcjczIDoCyeuU48cDQu0+GZs9O5bbN0zx7BrEcAgCTGQqQO
78hEs38+wd8XJypCTURzTiSvtapV6O6hEzdXOAl9omo84ZNIFo3zNpmf7cEV9hD71EIl8lRG8VDc
/PTSj8B+BjY5jjca+o0lyZH6sEAUqnNdv9gVavNpnwf5ldUMn8UNINxBy0RlhREMuUPEiML+8rEA
QfcLjGj3ut138EXkfssSbIE2IcfpYVb0v/gqPBCfgz3K4baX687/nQqkZeOA48eD5UvBSQTSGCqU
cUpq9WlP8L7Tz7fFT+oJ/4fxOGeLIcoefygG70SC8U4+Fgtq1wLgLJczEMpy2TTZypsTmJQyfmVe
AJfjhQWVA1p0MXM1EtYrrbezvHA9UyFn3tv+B/1g7l6B0EdCZqJfdSRBW8MP+nXzrX9Qlw6qb9Aw
QT5ow4eM92jTw57QN2xd3phfe+fnev1OzF3IafkoOs302nx7x3kcDJPC5NAAFqVcAmTamJm0wd3M
7DIeV4C6QUR0Nn+SrppzCNK74M6FZJNksay7YnpH2K9bSDuuRK1Je7RIQB51ILQtoq5ANwDiegXy
DhHeriNCzI8GGUEbspjDC3I1MEICfsy4bgc+997KKVzyGbHLMl4dUaG7X11nb3utUL6kr6zHPLqa
1cI8ed2gHBe1Lnymy6AvE1tGAENQS9yVqhBsUxyV4vB35vZfXFuGbL6hZsj0Ajv9JbgP7PuEnFKn
/7YSWiSJ1YnxPOTPZKAtqiwPxT1on4SZNsbGJAD24zVIlwcjMCGxuxAApnmvxgbAb4hiSudYJr3T
i8bWj+TtHXwtYlgqk2cvP20P3OhAQlKGTpBoedwP16NG0C//xlO4Ih1IcEoZhw1BohQPvLuFjmes
c50Zz3FBI2s9Z/K06RJvcwMpb724f7o03TuV/+RBgLlDe86VqRu6pVDL/je8DA7IQwYNVU+f0IgQ
O1+HclQp6xJ0hiMyAxpGVruoqX6DQdSy9zZ5Qqb2JcNwqq7Nr4Scphu+6J0ICqs0SJfg6pYe89bu
+EejIIcDgqSJdbyHnzssfeo+C/6UwViUaD9Ns0kqUgCYeQUDS3d2rFI+cbd8bsAfZyBJYKymFaT5
ngWzFEDS0/R+buKufOiLKgiKiBLGd6Z5pLLQ3EOJzLdbRh2wYCk5lXNzXrtup6F/J78+7OT107zp
BGGe9wb9AFFgePj45COSG/eSfMxLq/bpALc1cI0kUHbLME1DOyZjXAGbFzu31JRb6ekH5v3LZjpx
C9ZwObl2frzjb5WlXDsB86+QC8EH/N/onjIbbTBHzMeg5ikxASaqGXrA7xcqXvXetnJ2k5MyF3iR
cHD6twjA8QKRD8sAsyCzm0wQJqC176uqLbtMgRRKAs8XpQFcaWWPo5ge5XXh9xoaiJ2K54Ljcm2v
T8KUav234vyiy20dfWYXc2ZV3JE3lJJjAMIClwv1yBG6JOCfDEaXAES5oOP1zh+iU4g052lv1mrg
zNxNHwA7BRxJyek8yoowS4YhBBFv0EkBRZmybzjesJiNpcwpjxgKNvorf0z4+18tHIA2soA9uWo0
zRMMiPP3bQpJrc1STMvu1LIvf9LfPsvWsWfG9+R8Dzk3+Lhc3DeP+yOaOU5be25z2KHCQ/m9hCTs
C1vkhNqP/kNNNHzeZTG6HRZHPKGOY7zhvMkIHWX4alY7iEPykzal/dKJ6hyELiY6VHK+jNmZZgjS
gI79RVhIeG21GPcj1wVHFgIGeNamWbKAbcsNKs9n4rwI6SqRS69at4fFPoKAuLB3pKuXi0c0PVN8
nyvGMDQW6N6MHA/gAUOUUBBDdUG1kc0eyVEAcshUP5IKo3UYOuqxvTBideI8UvV5qvrdXFW9+67O
1SRiMlgAEkwpQViVNCWbYTfEpGEpuQGmfp6KC4BPmxJvnlnxSQcpfI3ZQ79rxo47JnkVVe2eQIU7
QOv6pGpYl/q5iEG7DNpO4zOfS0KnBJFdU34bmhvR1RL7gGxMlBr0OSz1A2kSoPUZp9C1HQSvZbUd
QJzfi5Hh+17ntICMZ/pFDZwKn5Hj7jYjSKA/eB9MCBRwuI8+FtQ5lNWo3EMj9swWArqlCy9XUmjF
fhZaggKLAZnbVjh2uGfMZXuAt9fgEdRNei1VxLI4XeRQIqjAclaKzewO7bWV/UOlWabbtUKQqWol
66Weiz3A+yk48t/UqRpv+lTiL8F2EcE8BC1XnBENbGggyXjU3n1F4nLOtjSLuywQ7rky7NxOLx85
e0RwQymD9s9UotjqHS7UMOIzEQRCzFll5p9F5NM794FOTvgYidm4EWmsx9nHmOKls0NY5hHYncs4
l2aZMQvxbldESjTWMICV6qTA2RrAn4c9p0jpwPrXjduKW1voin2w0u/H9STU6TRobvsGCEWa18XN
/txnJ1wGYYvEG+gWpYh8pRXotOzH4e1SyLL1pB0LG59ISRkbkI9QqLHZglkHQqKysfvZ9aiFNtYc
g/bNWDDT71uNa4wV4X8bnY5FCz4kPx9tznzp4SsNNdYW+89K5dM1iyus97pQTI0gj0Zb8AMEN96S
SlFCqj/uC90gjZpML79z3HAqKQpe2Knxv6flCAW2wh56CfSt/iK3y2Cmvs/nViBk++PSPMERcIna
+CJ/7c3Ir3BVncDs3+JNOohRTF/GlqKbEMjkyGeX7rxCwSabic5Q/GIMV8XGDxm6LZ6CfRJj2y4m
ZrchrU/2yzba5k5N9QP8Pm9L0kH0towNmoSm5quMsuKJIt6ePz38q3+DwiGW9uiCY4B2ga8AvBz8
pXY1LvV3C7B51VEUXmESs4Zoi3qb3u4niOSawix0E3KJzZOczE/oqeSfqRJQlEeQwvMI2lj3yJ+Z
+v/6Ilhip/bL2tUuJtZfFzJA9AU943XmdPbgz6f92iKe/WuHJdlD5TpERuZqYta9QCzqZyZ3Xjqi
wdkKGMN0BE6uhTSzsqg+WBvLEQOPsD9lAs1o9ghHkqAnRjx36Sk99Yp4wsOVxX2XKT5gF8tmhlGS
2+DZJvsk7WDy7EtZektZTkcrmn1saaeaCwSgTC/ysVxx4IFWGh13iADJqgHlXmLmgiFPNSay7J6m
Ku2Bjl25goD1Es3OzaUhgG9k2lM5ytJ6pcvDQTg3y5iA3iohWqhVEWvonaBHx+9E2YEiSXd/0LS+
DQ9CIANgA1LTUHsMFqKsePlQxq8t/G+cGYzmyRXe/jw4SB3Ec2e+4XFR0iRioA0zasrFqXqoFnH/
Xe9KgCjsL/P9YLD208/6W2rZUYqQQllQ1myPUyyz2Lo/JynUkJtDHYeZZjypx8PSY3kT6k47pByV
/+qX1hE4TG9pA4BRkWXP+Q7DG89KHQSd/UVdDsMqSib05iziidl/tDifj3LtLZDumI7mgo73LI4L
Ks7gH8XcJdKoDexvE/bCCeUHKkKwaxberTWLH4/gm9BXYu6Xk7Zbi2tyZR1NRahnBmRkPczhs7us
5Zn9nsp7LcqdWzW+RBz2gYvPSCtkoSs79Ck/m+7ZCBMMuCWUNDdp9w1A0mH/Oh00JfWjaTDiUj6f
jH25eOm/QqSN5qV29Dd3TD2+VR6XngHj5xl3BXn827xH44M/dv3AJPHz6IPnRTCtH+ckWxc1b7WW
IhJnORSANH4Gs9wurEgJTqBzpzAdFZ0y5wIlkKBZKmEXbmaqY28LK3HEOpywSHa4fDPfrgCS9udR
bON0IfUMOj/zEEb3+nh9q1YpYIIWRtbhpkrpdyknhIZbJb5EsPdKwmyyacnEK7RBxv7vlAj4h2Ja
RVhSk0lSGZuD5clie9C54BG1VqwjMhfCRmdKb9gibi+YLMJpyrKOdRGA4btwIyr4G9C5zKNM0QOM
PzVOX5nWkUglRJBSWiFNuLnzCmQWYPW3wdbWJshP6XrNhbEjgd/DCUskbRLgn9P9AA/RAAbJjMMF
0CFdGhbJ0T0cTYKTawfosVel8T6YqKYyzAJz7l6to54YHOLki7f/CfqpnPpF10vMkaFyEG8HyWLi
gq2gSv5bnbe62F+qrpng/PITx5h/LV3sOoGnX6q1lNSFxAtMuhkHcnndTzkUgI117+0mFxbzw1W4
LTCpPpNh2LJEkBATy10Q+Y3cKKL9cIJR7It1H8dnsDuOguOduMVauiaHnMB7WtEIPwRHcC3rId4i
jy4zGHpezg8t6mV0vB+7KJ6UhkOeDwWj9QF496/eRKtwAdDlMjxp24HSWxsVRgvWGeKcaADnnF5e
D+7Hh8WEye0AAnbZtyUSiE1oLnxv32zBZgbOACuPRqdQWX4mex5d6/pN47pr0Xk9pU1tGOhJDmCg
b1X6IfxMHslzhw2WYGgWleI6p2BiNtx09UY0+3mFHcnSEwj4hO69En9CrL0/RSeAdWZ4kmQG5X4f
zP1BoKCpxzLAum2PcbKVsb0UPrLxFO1ysryF7kl5R2siztDhql8FUjQ5LzLTU5C9/n3dQgqvvC5d
GcVqmjPoLOhWn4UhPPPs2NXD1N1JZTaxKwpbKplWRjQfK3iwzF3QiU1GIskwLtL3RCTG0WIs4UMf
0Fxkvaxwu2ireDXv8Z2vApgS7rnbsIqQDJPGiKXlDXCTFscfLDhppkfETD8gQCfZkkvmlWlQ1RIX
ujKsUYSc9/SfdXNuBe54mGL/APqmYCnh4r6rtoEdNioh0MBL0wPWnF9KyJ6szFmuNpK1u1Eo5BO6
v+udw75upoZL3198K5xZ8KfB8XXovdIahe4gTRM/4vInpqomLDg1CInI6XNSkJOt77G+HLKhK5ux
eD93HK+doWM0hRVIcSpWMiRYcRONtNezRj3aM1MeBPFrX/NW0icj04PG70GQM7YSZGOoY3z/I/eN
WJR44lzjmZx0otc9fImb9Xmm1nlE7AzDvt209y8zVL6o+AXSTmjR3TOWEiyDBsGw5T+fqRmZXS8x
E7bnKFor5HO0glFeQF0sE2aCn8k51FjAIa13M8eLazVc8OqjQfxtPe6x4Hg9Bz7EKeYxK2xkAsmB
wneNX24b7/+EmSPfaflhUi5QPBwBgxhWjKsCVqZOl+cCHTDlRO/MXLxl4uoF+zqpvYfiyk+FLud0
OxHOUgPe29zhAvsTov0kFFXDGslrtOrS7+a46xrNbB83ZBlptHk8J6g/LusuXdftU7tF2wDqUguS
DgupW1WngqqfZ8+VAqEeNDVo/MqphZeyUAiuxG3+zesT7DpnFa/q4VNnBjoqU/DFfx+1n6hb/qBg
7ftsh/8rirH60IehF8ighNHqvju4ADIpH36vXP9XPkdP1EAlLYnVvsBlKyXivolMd7OFH8FvQzHE
4M8DqgBZ+1TH2EpFeQeF/Ks2iY0kQTJWCTeld8UGrdhbXrXOgPXgwbIwbDPUUkSrPrKDJs27E2/u
07XW3AAIjVH/atKs0aGpTjPm+HZQXBHsYBCsE4EVW7c2N/iqtTJmdSr+Jcflohkzp12Ho8D9KU0b
c+FgBcLdxKZFQ105ruwgiOkW+N8q92B37oPVQoa7CWVFxWSYrJQ4klgRDvfVG5d7cvzogk11rivG
2nmvseWOvTfU7bwC7ywNYoYkcSTO0AebE/VPIG4VStC+7eotrnkwq5jHySCqcWZ8PYKZlmYC5Ekz
G/SxTgR2NBZuPdUHkRIJ8sgpJAGvVly8M/kqnDZy237MZIEvzlYjduiBYVMzMmqV+gOidT1AO0ww
voUgrCEsHHzT0tM0RZ6J0kaMm7mI6xLYUVBSGPtgO0+/WnaK486NB0D2XhuBGiEQpx0d/yeLjF7E
Ywul5f4txKOyVAFxfKo6ZrDmDUKEw/xJYwrcLNmO8leyUKDVn7MTv4CQqmVwsTLJd11eBrvCBoEy
FfB0+w49LJT4VVtb6tBTTz8LQi7wpA1kHzJktEUEOQet+i2atUM7z7uGmvbhQHtZkT3WHrUy2erj
rwnxR9F8lNWy+BVXlBcnOHu/+uMOg+zY6tkAr6gRWe+D/EVPOgRQpUuzDTGTWD8F3QPvpAAxg9ZZ
UfFzPeWOpmdj1n+QaGIhCLzX7ovfsvKdnNFOzB9VZRRQUVfMjjHiNYoIJdXt9BfIRovdStwEyHZw
wZxuOIeVN9Fnr3kMr/PHLUEmLcjYDKb3lrMIllO1+PS6wNZ5a1GNi1aAaDzY48UXTk3CsyhWpTdd
fy7QvMGzp/dULxRLa8zMdcVtINHHu8Tgx6DOuXQtZNMGBp3CppFcSbOZ6rIIjDkGnFRTUTOUzEfZ
ze6icYQX6veDHaf9FMBbSxpZjhh9YX+A4Xh2ya7NsFbXRb1VxhVGyQznmoh72e0LfJwO5ktGz+4m
OvD8UQLCGI2ShgfhWgThY3uNZMU5CM96rrPVE0cvigikkV7WJH7XEoHUeF6gp9UHgBBg5bl/VCtd
lesAeEdfx7K3L0w7BREg8rtAWDMfM93eUzlvYlETBr1V+cFqpRmjYsvcEOVCW9Xc1iI5B6f2ywCf
RqM+A1qarSITmkjg+Zo92RS9Tsp3k1bl4BjaPdNKCcpUmUVrFzgO0FEhyZuOmMuGV2jZPkt1E4ng
Q5kU0DYSuUN1xlvznu0N079up2gZEu/wq5QFQY29Q2pkqVjwAk7X8cXd2p4rZ/WeBmMAqHUwui9e
enNH9mhxW+Ft3/nVan8GI0wTSPkl9VWIvz18/bHaBVPiBZpsj9nWifrPE3ffWikx3h8yZkX6M1dU
5srF9QpszS5Jpd6doreVVVmrGMzXYfI3coQ9iTjMe/vo+Aa4Bushbw8GjoogWjuwr3P1HEJJy8e0
HkW8vIT6MJsPtt+lPzMubwQSTSdq0y4y8fGTtVoZPGk0C8LsQ8paRBIJ7TaeFkHA4jjO2Nr+PlmB
SXXHMtJfqBdjuEAlCElHkgWPdFmxfukxFqKFnYbkf5EvSAAbd8nPl8kqt46rJyJJvHTSwINQ2CYu
eiOdzn/F/UP46OymC/dlpZ7J1PRDNyzVxvSpMMkrjFLB9GBKtDOh3IWAI8SJ3nbFF3E80Ep0Z4rK
C8UFXVmnHBaQGF524ynFjm58Fmc3NEL8C1poy20a/O041CWfANN56MQqh+xox9x28vLUhdJmkE/6
AiVJYRl7Ku9wI93wmldsSJhnOJD2n2vRB+mAs2qvU4uqSJikCfWmLHmSdyx2jhDIAazHojUayItr
12lNjCu+enSsm3tC9+33wMzLjHNypPe1vbg4RuQqsJIhqA/xe8r4d/ht/LB2T0HFIaOlgRuIoMWK
EEoTyMuqtXKT4iR9nurYUIuYJP3H6cXXx1u1lLjEp7lZh3DS14xVB/+m/w4WFYRdCBiXli4FXbz1
9blkc38OEWBn7DJNf1G6KC563+Pncf30eL9+VGYWML3vRZxRqblNigaay+jYXv5W0SOhYbdmxLKi
OALS33iwLiQAdzVsvxRVO5IgyGBgyopanCxj7saRILMBprKIwvCOwLL0YFqU8vGOUpERqpqe9Uvu
GmcvCDnWzwm0+0MV9L4YEWm+0zMzWpzdw7XL07o3TNSpL3PiKnlNCR56j8VETEEfolcfywBknQtY
j/b5tdhPGZYlYMLB3RQ0kp68zs/0oUbwPcyXT6znz45nMukn86dSEQGb7eou2cDLLhTwfe6f3SVx
gMrgx83LNlGgCzkY/IrcfFY+2iSiNwIJhTKZ6yQoWUHce70EU2FmznNxZL+BLJJH19t02ktgOS1K
FsgN42Qf4D5nBmT0fqRqPKUvDL9+2BSzFqKk/25+2iWA2Vxbw20OJ4ZwJPCl8zCLwk6hgSytAmDh
MffS4sWiP00ySifAC0a/KHsNtWVL/NC04cPFH4sfaNnIscQiBNLJM7TR92bPGFWPo54Rz/WGeBw/
LNINO6HKCuHDdKS0hjk3wrdzjXO/EesyChtdRhbh54+PJ0a3mPFjX/HZunsduE3lmMnd6hBxj//8
QwYGu2qriv3vqFWvQhZs9UI3Y9U21AtzxjFFb7/ubzOqV/quZ8qhP9oFGkbE26nMy36KUMzm3khc
ym40KT38ynasKcpB0by/UDT3AnwDR9+BvEBQPUpjNyNoM7+Y2yOl2LHGfjZAPXBItHtb/WC+7ir3
JEenE2gLML1MziTpaLs/03D34XJz5QI/S1fhK7jPabJABVAnK9S+hszxKeWt0ORQJVTO0kqMO2aP
8ywih/3RH/d8dQcfCT3yeeyjD4PU3vchlHokMO4/jWW+zpQHNR5iep+4eBspOsMLmaaSz5qvQ4TX
O+tf0CrZEo4fYRJDPjkqXJXsPrs4YJYisMknviW/SenW43wDUtM8Rp81rl94u7snbkaPtYy9bXse
B0UTSw07Qz6LBuDd2PIzk2NkmyQMeqtp9inu8t8KIQtPtT7/8uWllQWN8bzr4DNKmOcL+hA6nRgq
vH34YotBU9Cko0TxTyYQyJdzxSJgQgW8ve1hgMY0a590hlMYEuOfFYGAEgzOFIwGOy28mWiz7D0O
AJZLeiHDHvAOTuhOYvfTyQzSeLwGRb15hj5UWeHcjL/uACdlGDPkGp5WbSXFs0p+Ja16YJjARAbx
5yG/mETpRXSte9YIHUc1UjPBEpDzsZ5sYNBR5ojoXSj+899l9pf934Rs9XTrtwPkpbhxTmS0lCr4
YO/rIsbz1Hw3lYSLvwXQ6lemWIHlDo4ISKPAFkwH8mPfKeSZXnyYsaY0mZsOdxUQ8ZKKqYeaEriG
mZVGpzUz3j2SdkAcTgyBNzHwYWrddtK4u8XGyhRLsUGtXUq/gZq7ItcuRAZTvD97g/c5ZPLVMX1z
halZltrz7mK9OMuY7A3bTgHD2inEFbqVfoWbr0oJdxX0WdHtPBhJqIrqBN82/YCDeU7q2Tn76i3v
9LhThSvt1eu2u7ORtCLR7jzQsz4/UQSokLX3Cs/4COrr8EmBWPlRnXJMQhknLUwo+U5UiWo2NJ/B
gYfYii83+2QYG37JTVy4GpvObVa8U7bDUluCaYAkrMAfP2UAbXQ6eXnOV+cumJ5eyMoJ4DJp5YOj
xTL7US/lEAuhg/IXJCMcjhzY5qDCcLfJshAAoLZxeY+VQiPVXuiv6Vb472pxtk1PFzT1ENUfI2dI
wm30f7fSRuhwnaK/aRj/hWJou8t8rQkGZcrq2a8rEZaMCr/eXaSHLNRUTw7Kamp2i7TEBlDrSYpW
FkaZpkt9JjGTj4P3faEfEqnIE/EXEpaKBxBG8kjjfgG6S3kkYFbcZhTR/dh95d217r+S5uh0S3xX
5KfOqWH3PEyKjfHzfKw/YA2tw9WdHzZ4NZBcQv4f4IVXKYlJ5F58s/ZSVmuMHfXguL9cFfm7bWTN
K+hjVcd+P0I0RlYJNr2zSa+MClNPeKB2td3CEp7vuygPvgfV4ntzgIhzqv8/ZlsRpg1cNgEXoWHO
8qQ24S6ej++N8acIrOKF3ifAQQRXe4Y5FYjmNEX2T4sz54R4OK2xZaQZgoCh4MQu0MrAVc4aS/RD
qKxceOz1FILX4jFyNsVojQdODJEAaQ9Jukcq+OigNBcU659bV9FQkW5R4ZqNhZRZREE3zyZISUik
Qrj6pMPmIYsutvHTzdefalDLxlOLn2Zqyx32/H7bazQg6QZDAAsM594tab1jWtTfzXlzl+wcrgHo
VcixkRXVdD67ASN6nytoeizGTO4mm7uAesDU080CX4uhhSVZJDLjHTuAiNUvt4wBgq5QsdPcmm8g
2Mw+VWebFDAEVehtevKVpo+ua9ZVHO99piXIoke8/ZlIVAWTws2PKB0GiR8L0i3g2ZpqjndzaH4e
pi1yorpVsK+eEO8/cKCEamOdOpuCD/n8PZGCntg8SuYJ8ArumTvUpzpq1hmK7K2X4CvEuwE8Obg+
ILQyv95HA/iz19fZhFfiWxUb763wzoUoc9lTrvUnUrAEzgZFSDyPLQb+VvRJtVB0Cbp1ewFC6YDi
jWVDAVmBqs2K5Ir/E2iANdkN5Ta7jjq7PfpU/S3TAPxBozo7m0EpJ/F6pnxI2cwoxJIJdEKt6E2z
gcu/AG7RbQqWmmfkzTD7wpXyKw1um+obVwsHyqbxLMZhU6RL5va5Lq7AwUai+tDLqQ7PPy7uk07f
LMFeT/Uww6S1v+NjqXq8+PO1nupHd3kWfbyeKA5xk+U7DgoK8jxhn5Fow3XIb5oPMwbhq2AA8sjp
1fHj3hFjCLElF+Jd0UHb1qC9VvKZmibR855sPmkAy+WDfWKZDb1VAXRigYYUYEtUuzJATEMae7SB
nfr0/dwQRqD/NCUjuBsbAuxWhuiJsW9Bl5mZBPhUfqi/8CShCjUVFrZrtMBpIffKX9sRSnXdRrfV
yla4+V7ml83/ZiA7JG1R1x88B+IgqtkycGZ32TBgG6pWMtyya4gXItYKeMlaOmegkjqnVvwjHiNP
TeUzSoluL5NU7TzvysKLXsE/LKR4kqMUr3toGhcC7LfN9rN1PsElqD7rCdspbTyMiseuPzfhaamq
47b0wdoBlaD4HhW4G9PIt8bG2xbjEi/A7VPqJnP6XfH5PJhGpksH2u6cdCypz9JJf0Y0CK1y8i9+
RWjrvpw4dM2AxwjM+ERzt7RHc/vHyNuRJdaNemvH88N0xz/EusHpqchV9RpdY85PYUIFONirdRAL
s8s39tTC1Icu0hsf6Lo4cP0Azu/nEHwYbcBv/4rfVb79ID2Nu0S7qNnrswTf+HOIWAkrHIX/fxNF
+sWAQlzJHUnCMZmzRRPjcm+dGE9njcplCquf0bFTHpoOFXZ24LYwVkkByHzKvH6BA7YXrPPM/SbA
M9Bh8hEb/2JIHJ+CAgDCkPgiPacynnomVxFsI7XfR2Dp5cwZqi8A6pWKak4Op4FLYlYfWpf3QLzr
37IxiMnPheAEqG6ccL7WJc4BUMaNFitdFw5ig/cjG99CSpLlaRvMNzSATfvCnT9mD+xqTxCR9A51
WWUJERHBhSo9VY6IhUWN+4NkA7ob8DLZzT3M34oyWRfUmdBajogp1s7zYauOmrnrpAzNYoXEdQOk
FvIFWmgfIEn8t077DPbs+8Ho0bZRadSaFnZU8ksB6N05C932XQYzts9rSqiewbFV6kqQW1CoZ8kS
A9RtwxxfWf2n2oLErNDjBou2SWbBzpTrxxKy/jXpjsrxSZCmlAxp6qo4IO1m8VO1YjMMsHVf5T8c
s9tX+sK7CJju3QJR8PcLXHY+cCHecf76cAZLn2UoQ0DPgu69vy5Ll/eKyqgBur0wsUPXucxUcAaX
KJwpDmGkLemaTAcUtq85lA50x9vGPqhyFgQEzY4qlbgYaZCkJEHVRK5W5WlfnsGRveivEBSaVZN+
0tSTQiNd/k0utTWMcMGeGl6wDouABKlS3jUCwHr1WXWWIxv28CWjI0znrhtGVaZyUVmBINPB7+M8
pR0o5/GY1ZDLlD+lJ4t05BzZ9V/jJmxWcebeIZFjADLikkKfBu0rEfPU8GNObVEzHKUfAh3CtAmr
rHCVqcgpvZ51+gtDlmOYngXgFPsc6OnWL54Ibiorag3hp0aJVm7J8KGN+eYukij9sxSU/AyGLjmy
mLcevHN7FYt5cdPNFV8LB43xMPOQaYqMGOKj0SAdfKWTMgoV3C1Y7jrF3609DcLi10UJEJC1p2M+
Pb2dry5qRu7xhxRf4hmRpdX9uFHoTp9SXs4i5YCKveE2dtjJwODsixK1Kq2v1gGOkXMaQDAswneL
wMx+DFS0hJ6QrEb9pH13py9rqKAOSUkH6gDPSyMA6qMZK+FektpGdEfUjqiNBiBCYM8o12M88wYF
4PjYNLqepGObfmsa11BfwJvyPS1JioLtmTIVmxJ0QMVYf5BkewGOTiFqLRTSN9zyJ2skIQDowSeN
bEEs4cBt6Mt6wlHUZyEF/ybrp4ocFeZyT1tgeyTyy8xmT2weUjLNM8LUjNrIKR0YfhVi3NQtoCAg
33PqcaSs2hPgsCkeoOx1KCUU2RuFm8MVIy+s+DlK+WtUoKUBu9B2IswCgjkqYAqRIsSC/DNOUSbr
/opJgyGechVstNSL8FKikajIR8pJ437zE3rXiuHxbXEb0k9qkwV1hkaTNZxJzoDBDPrhqFmcNO8M
3G+R7VjjiGHNHDiQDu7tPo+ZGHXgA0XmErJ0gAwMoRFDcfrGVuewhfebDtgFUKwD2UaJAxEX47Cc
zacYAchXdjZ2c6XszJ8h0mInrnCE9Ujt6lnYNDlomev7C236oix+i8wYdhZ73A3W89LoI54M8OBA
fKAo6mURFPKL1YMUYXMDm6B6X71pRJtv0oRn5si6NtGROAPsvmWlNVzmfmmQBz3uoIspdPDwr6Zu
CZasoTqOv4Z8GR/eS3QCbYFKtNz4pZcecP4748s/QNQncbTczgPNRYx2hK6YlaeR5GrTLg56f1W3
5Qq25cEPCnnDW47hehrvZ4/D/W2SJ5eBIQeXELpffKvJ6VZaEV056FmVoC4rSscEZ6vB29SYkja+
FaD4C9dYjXCeJnCfeAwFKKFsLlWq+3JopNJEgzIPP29DaL72kVpceNHv1Jq8V8mzVi03jYS5zRly
zz8wrb+V5a/mQlgt4u41TEdyJghu3HzQvihTD63ibonU4BfayzKtJVWn6YjaqzcKLiFmNT+PSD0Z
QviqQXan8Ppfa/01pG1QFZ8jdKaU08EszQfW7KMRr2p/TuqyJqcgSPy2+IB+nSOiGIbHqwNmSldn
cP7TxgG2dfe/Hs+3twyu50TB9Gu1spzM8iSopV+5924eDEBE3k5X2oOfMzUkoUZBOOlUvAqKuY6Z
7lWPGOOklLHp16dMDEqFTXYhT4eS+HCYfyCCBbFCwrRxxCDhphIWSjKwfKLeqjhC6fqyXKuKbrRL
i1GwClI1BtRs5pZ1jaRAcMLoRFwVCweSSM5D+EMp6NsdHFd52V+248BIBDFApZdbZ9JAyy09xj8G
b68qw+Tn3lFEdinR/bGcQNU5YPCNh82mUTQOp1UgfmAJH9xjs4IIYzrXKaPqMAMgsYa9qUE/uEeW
DVdBO6gO6uVoBOgVQcy8a8NmjFW2aQauw8qSo5oiURhkDVLMogUo/qAvEkx3npaQ3CshKTRvjRmz
Qr3li+n4sPskPXZOe3k0AQoyPd/b6MEcqyCMrx7mLOlDl4jnqvA2cpRVjzLLeZrUDOxiEKd2CBry
M8uOBRjQuVl9CesY/VE56UGKlAT83izy59SIrFbRLOy/Xf8NDAo/8ubwOr4VbNxPQudl+D2x+miy
WHQti+aT4Aaku4mLPoXUNeMHosK+ZGCQh4rNIjZZ9ziKbSzcl5m720SbbLhxtqUX7ihEDldwzCPm
XSHA+yGZC2y+RbLvht9orckpIMRz1f4PQizbFJqKUoa8cTQehTDen5mYibya8H4S+KytmH8KUVUD
bplWfk3Dat4jgFLriW9CgFd7egbIG8iohgaGD7KGrSWsfvvL+se5ewndynnUpqFtacdQih0qYIB5
abua6V6BTPWpByR1AUEyOHN7IRG5XvXQlKPzxjETa5PIy5fcR32WRFvvl5gF++ndCPRc/CDF9g45
GamvmTa9GGu/eqN3zvai7+V90D+jPZvZfAfc8FjTAAJ8hetx8NHA0FqRp0bvywQtEvJG2Bgs5p86
cD6CLxHCDNYR0uzqsSe1Fuwra6zVgYBKKybtTUgB4BgIcaTZMEcD32OF5SBT5MJ/XlATmyOKF2Fj
v7TNxTDzUzdfhkNqVwlzwWOTjrEfx+TOLMLIrvxy9iJDJGv5pUBFebwc29kNg11kS5v0NuPa6Iw3
5lplm0mSTK5QfsZhgO2A5MdexhNZu2d7eZ+Q/K3ho8wlFc7guQ3COE4VO0wPmZBYiHppMK+NbhWu
OcrRVHWGbm7QSGeEnLPXJgK0SFE30Sa6m8wIGX29SWghL5jJdjHfr6ys83IKZbUY9m/22gPv3Ess
2XQALsRHf+HaI23h/IMLcbG+s0+uB3yr4qKZ5qPCkihb3JbQbN8+FOUEkeo6PYgSUe/Jqe6tebCn
dzdQuuQfYh2digA8EKgYRGc6l/I9hQKvZo6cpBZUKrwsJjz/5tmP+/O1EcVNo+lQ+wAYG9HUiHwa
Zm5XN5O2MpxmW/wnr88RigpweWLpBS3XLLo935qprsuHwahCrfDx2WCuufiTCwYu7Eg4C79UWFx/
FA0CuMK3fluEHJik8mIJNb9BU83/wJoVArsDtlx6m1Q6Umcjf14ELOq5BZZa+nacPJi87/uzYzdS
4jbL0JyW5NXdNAnre4ZAU3z+0z0c2W7p2YFDUmfbhfqt2euXjtZJsHkvN6VWzFqjs7HtxDFoRjCk
7goocD7MaNyvJUm5QbrUTlsylcYDLUzvdGK3lq4Qzaj8uB7EfGs8TTHu0aLuQbIGA92AzDlIdddy
QHrvlhxg5PRYqUdae7XL+nIDXkQsZDW1B0rZGX9r5mVsxZMzTWjtq7gY1AgdjNzRaeGpCw8vN+62
Vu8saV65FjoTOVzswuphnwJ6zQNRu/QqVkZ1mNaqggl1TjPFZFH4xL6yEZRLLk99wB1vFXhhHg1I
BfmLUloX0dTE3Rd5J3cBk3NG2svmNAlaMVnk26ycJrNUsQtgbOVV2oQ7OPOkr0E4Za/XE/uOQR4O
co6leT2SPZJsYf2D2vOUnT/qEsuD8fsFDaknVFC6/F3ZRs7kHD9Gl+NHbydf3+MqLNp/DkuNSZ6p
51/lUKAUhYsxinQ9xubjgpwO4zGSBUcj6ZeIlirB+A0tQOpdExkmxe6cNpcgdtf+Pf2ezwd9mGsu
F1BIsEv43xUrsq67QyxeH7Erv2MPNKMcbyAcugNS5dQiFi04r5jFs0Mmv4QppVBFaewwcrqwLLJE
ZyBqVPxuWn8gNEhpVd5N6cjUdRWGEC+X+PAyyxEV8ONqd5HEbPUfU3QiyOcypWR2ilSaZxm9gJce
NjR9qUx6VcaLNHRBb6tNWh/HQGQwDykYJe+PnmbrGDUu+XiaBsuAh06xadBCQO4PqF8QvuQsbEL9
oe/ZE4k2hcXWN6aU6y3v8hJHlkpYIC6lHN5LFJA9DZuajw//8yTTwCBQbQzbtfrA4TPQX5l+wj0q
EFE7G01YEPULp2XqR2ZAIkrGwuQuI1QpdoSvwSSTT+yANhtDg1JNu2a+Pk+rMNtS53Df9lPDP03P
KFMvm34OyV9GmCltbFGRHYR4PWkCZCbLcFme2T4hZWe9fX6YAyhD6McnEVPEJNwhBCazi+sxyTai
fGkkjk9J9HU8T4vvDrZ2A7P1zsgQGPcaRAjbCq5IJivTPGVMboUJasfLKroHZBOrJ2PSMWoOHWid
XF/LvTw786ZWcj6eLwg5SwIiyl+4u+Kc1cCZ8XvPw5x5JDbx1dyixTHlnU0bGlXrUrdjCgRE9FNA
nk4p1ziFLK1odldIMA/LEVXzYhi6kNfO7kn+6y75TEb1rP5e1n0YoroCQ1BIQ3tX5mGLRhBNqD2f
kNiY5qJcB+jZax+faq7lav2WLMm6zt2A4kdADyGJW6jelpLIWnzUt6N0odKD+tvfDcSoFtV1q5mf
I+GGGBKkWXy8r5ag0apvVoDJaA9AHX2CEJK+oLPIIGIcD1yEcfo66PNtEekA1BBKH44tfqNi8BcT
qwFiDQpplzU7ZXmZkYqvTBM9jdWxpg9XWA4kLiTUZNJapW8IXUGMRzAKbdfxDhwzpOGzdwJMgw1b
BAoZnUTWROqhadwXI/a1Ug3Nkj8LS8S0skzZ9t23sFn9r9HTfZwd3hVaX5OZj+9QlLMRBrwYAwHn
pqJ2lH5Z/B+ie/iYe6vVwgOUzD1iWHO75qUAn5/2AoCeiehALQpTVB9ng/KlQCPm8XE7s9QX7YLu
5EYGZjvY1iXLXUSs8a56nmYgMNLSk7Wx8z56G3c6s+Ji+tkHnbjbme90QuxqWPsD2q+Q8SkCEx3L
XDHMhbPJRFsAeJ1stWSJxeq349+4rl/q6YUNvBU5XMzWYFPSmUoQKLGgvBrFE5LPkQ9Je9bn6i+z
tUXA5tBi4l5bCLkuv4hqE6Xyu8xWHfBxJKrUPwzhGL3ggBZM0qZdZBcgyTFG9LNUfqPdZHOBUIDt
xW7DGUzmX7B/sbzDhKhXb+J18REwmZcv/Q0vTga4/BZm7jIpvBXuz6LTZzZJxaurzHXwzYHzwwC1
6UbtJzllkhRelytX8ZRw+CnfkoenR/nFZzRkZoWT1xF7/3VrnSb6cVJvvXCpugiOS5uB7KYhZipS
ADCnTvMM6sM2aL7X6nKXMfnXbkT6n5KxOi6JnlI8wXyTyABTKx/BHjWaV9tKm/iqeLRLAJ6YBdtJ
ma464UJbXSSEHkwgH3DWEJMFzDo+IcXX5e7GyLSLSK21zXTCsRuJSYllCC6HSfrAQtCxV4FR/xNH
ME8a1bWlcssvzOKkJsFce2laZKIUxznyQsVDbBhqj2F/qwfiRrx1Jhxnkywm7HJC4njPLAi/DYd7
mSc2a1tnZsE5G0ayjdLJZmRuFWi3HrW0hUy+34317wEbSuJLRTXJt4VvEBuD+qFSPIE5cHcWE5qf
IOKO2473gicL7gYgj36HSm+tm1znCuliRR/kfU0Pk917Tg9ttaC/Q+OHmq6BlbSCuMnKpUd+VISa
GHmu+Js9f1gexUXgSTwmMBicpT1CjOr7KuqLHmkF9T2YV6NjTIdzxpgVGWLfnSlYMtrPxqRhW5TC
Q3Erg0IjG1SqM3mLX7jlhefeUO8jiKj5ryR8N7M/XUj+pSr3HfODKJ8xrDu3l8nagzTb5/QnjdrO
PWIpbKnZrS4JeskH02uXvTgcnkFl885H2zir5VaMeP/d3oJ1S/MMdjgEeRTnDXhc8h9ek9TH84PV
zlIyHGnPOY+dUKk+VtTPVi0mursQXf5Ad0KacTpkc2x2l90WJ0m3ZJsZPBrOd/pJs+EEG8FpoBEo
3CF2qR1ZNInn/+dXjrX0vkmJQQKhb/9t7ActD0NfHI2UgClwG45D2O3BD0+zbBujRQzmpXn+xk5r
IGDpG8T/nhGCW/P3bDnOOVtQ6jvPCFCKOXKRKIZPhSkZYsyOh5azxxJmcqcjbKNOPfLEXst1kloN
gv8v1uXSainA+Af48QMm7Ttq4WVbPoZwrpP+CVes6FK0K1cfXyDxN1ClvFOY4QdGUO62gU2+lHVC
p3CDkdvO5AzrcZvRewgPixDWUjul8KGxiHYqDIVWsyKlm4G1jPvm9FocxrriMaLlazSxv6jzNHgZ
s1axPVH1LJRN6jLq62JHf0+3HH2N0rc4ebPx+Az/PVwfoEJVIhk8LMfQiFey7+vlemfrNDoVpIXQ
SfdUtTjcaw39atODAhLRNxlHR6y2elxlbb2yuD1jlP6uZkI0XZIloCdirKCN/KTcxgwoxz2M0kvi
hbOWQHAnqcUNYA1dBP8B/SkzoA5CIfpe1YORV+3r/O//Gq0rntDR0DCiWueDFLNM6tyDmyBsIBEc
D9PPloDDBEmIsUd33IWuwqNdIjcEbBYwqqcAZ9d+1kQQrjVuDilO9R7mcNMMBx21ngZyWnKg42L6
zFs/gran7UB61JVqN4+6Ujbg1B+KQiGxuIkp1KDa5PN/VD6qAzDp2Bfpgs8GyYKn//kQ/XCjPt5i
FAGKodaQd9fv9WuXK6t5YjPx2u1oT5T5H75h3ZBj6KtKDKJpJVVZO3kTO4ZaxeX6B6FSwzESftMt
/7s/LBxvkOvVyeRcBG7QNgdXYGI7Tt1c/VqeimXaPrYLoL/lKdtfLJPqY625M+pJDbc6bPCpz6Bo
/hJhErgG94prr2Hi81ITMdwnh92ub5YpZu0N/GuaWYRYpGBIyhn/xNLAmJ7oEvMKzmIKVe1p5pLQ
vurAy/L3zL1btXUH3+7JzAMXrzDRfI9t8I9FqNJFIMoym7qRZ/6UJ7knfGe78rl9uuMFqH08l3Fz
PMUtQXbc0LXvN6USDcHXd3B6TW/gRbvsV/57YkYCBADUkcZJTlHSfm8+8S3wpdK0VcuIq2vzmOtc
JTumm1rW1Y5FehmW1Xif35G7IHMgchjb5sdIZtV/6T35Z/sgOCV8btAt2QYxsuf5zeGmFTD6pY8h
3etoZVCvzYL0r/ryumy7ahOUNG4q1HYEpv+A9OBiI0Kr4HmKNTUS2ON5jnzQFtZxgOUUxcxNLCsl
qfnXa7IcJRXn1c10m7eDQ1znBkBbEVAjwLEd/IfyTWUPlp9hhQ6n5c37v2HskynZc5aCdg6KSRNX
aYvKDz033ziYW5FLOdINdy3pOsGua+44STapkvGM6Njlz9HtkcU1pfopf/zx4HQet9W/Kzrln1Mr
AxePzBkfa/8cSXUtoZpLO6XUJ7IsvueT+Q98h7twb6dtHMfYbkPp0huSlwFbOwSGauHvTH7xDzMa
CDnwzOpPOGAtDNcAkquaQwoQvGNcXuLaBoEE7FyUJmrT+KfuBYKL4ErqLIDYagf3KTPqwe5RemeD
XJl5j0H2My2Q0IMtSNKN4IjEoFV00vRAHXu2KW+WfKKiZeQjccTSkXlDcCcCQuHa1AAJeAJILKF/
zq6rDqNfjmvSXx3q9nESkmabJI0IPjHDQcJp4zzAuBYYHwlsE5QDgcfRno/Lkqr8jsu1d6dwgQ9N
YCM64qE4Tplrc4G2ZNiRtMHG+C2yLed2y7kM77m6RafCN4gG3R6PmMA66/v8vhElKWQ66Efe/shF
tTUCujaHpqDIL6dBUB1412Ns9yZvoE8Hupy0ayeY9Y+m9L+N6DQw0ifgGF42XZ/8gUg86gpzyogR
1GhdrSCqeDqc/QiS/c6NrcFS/mikaRpeEYhSS+bo1ipZmxHdBhvXWs+8WFAZklT3n4FdbhGqJ0/d
mAvXcly7hwH4Fx6Az8PLlwDCSZGQ/4e4nMZTcui8SsYc8bMy/5Rdw+ihyl6FGP5L0Y+bfkyUOQ3D
aFhu32X/vHZcwiR5mvdgeUDHeUdoX3rnhXi2Sa+CyLNPF8vVZt677xhvx7PIqJm5g405BTaDvoxT
MGKRqwgfCac3TnJNLCJtAccXj/U/DVJEyiC9Tl05ImxnQoLBjLQz5Fnp4v/0K85N9w3N9NIh32eP
judQ/3TQhp5ov4pFLfpNQKny8oBpWToO6uqQvH7gxzWMWAHhxG0RvvhjSGUZqwbdTJQDlMF0HFVm
+t0irGm4r4xzOBWJl0jye1RLmo+aT2tJ4IRKU2N8Pcrqlq9WubWdJouaNG51iIRehkOviDKSykPi
3FfP43FqWg9qxMtpIyXj36orCKMythrgjD6oPigYvOcvLgtuaRoHlp7t6iwOMPX2rKsZuaQ54rRd
1dpZsJPtVGbFuSDuDBEIhH5mNq76fp4faB3+ibJJKwYmAaEMXyha2wJ0yvdUgcJcTz4kAsOqdLz+
dGKM71/coMjL5WzJICb/DJF58yMQSU4/33Tky7vu0tJ9oe4fpVIgyrKb5h/FMeuSBvAj1lLtX50T
AkzC0S8Hv6tBTIacv1qkvildsvJk7IIzfsvpja0hxhDLi/0kzUqf1JC1gjm7Ql2HawQNMPjp2k9C
Kc7JkTBDwppeK7bYhJW0wNHWmjFrF0QF7F9y735O6kUEjieoBdFbGf+fM62V/fIFeveTbhsf79fn
4IZehjkVUIy2EvuZoUp4rXgLSS+VdndXbJ9AzMj4J8F5QMRzyIjZKKVZ5DGSoOfX44y9o/bF7big
z0eiXHYY5M7xCfTczx+VaKDgaFEgDpplPnrvDXVyDpk3VGfHMaR3ZDDwJOZ/3QqKpkVAwrgMIKn+
62WbB5W26ViUbK5zVj4S7CrzILrUh6fyYaBQ02b7qEb4lM6rCC7IWNXLqBJd82Q7uqDn18IDl+Mi
BKPLi/91TUhoIZT1pAYuaAydLSlFC92O7wE5AH7L0JA6sp2sjGYwk6GaQfVURrzZNcFrSoq+vZ/X
4t3TSLQjOx12rJoSZbtex4iw54HfhK1iMMmc5Qx4DZ49OHZOvejgnNsTrbdpwlMC6pwXHQ+Wd4Vg
bbNIERPgIJ9O/q2QkhC++aYNcwbNIzhC93lB2G9srj96ydyEN5E6OBm64lVWpDG81dpcWhZQk99E
NqgagToeOMczAVyjJT7QPBm7lMKnn9eXLG56PnPdm7/akyE6mkbmKJq5cMt7nj91Xz7I/71eo7nC
n5BCoLV5YTyCuUXoiVFzpM9fH8CZLrnJZGU4xUw8wc0EH/dtgT5nJCKmRLHWhRnTaW74FZMx6UIg
aimrAJppV8xjHlhT1YUzUu9GoyH21fzPgQcrl2Xp4UlU4yoEKuch1QN5WmK5OlZuHeLGMeSYs4f7
5Laufv4+Lnk2jcPo0uw8J06tcnwSz4qeIIx9JOVITzh5hppxSGwWG58kQk054WuUxqzQdGMWTr43
KPG40NGvb8WZ1EAUhLhyVL4nlPpe49EjN67Sz2LauOTtnyUjS61npK8pMIK3L1DXSK/0aLceE26l
JFhdvO6NJZ2DKQA+oKyAxz0j4LI9MRglZ7nb8QY0t6fg1NEtdihPfUnUMhfNF/aw/rxXBXLq8irS
9sbdcZdv5uTcoVtiLTYyU0dG0PwY7RxCz+dxAF9457O9ekS2u0lC8APuQuL5RJp96yFvrPdj15zh
8vjS0teTwmwTgPV4SzK2cA6n6EpBOAJhz4OBOqvCZXFHTbiQFaTEiMbu3+scSjn7ejI4EPmOkBi2
qBP4vI5y6tn4EDEPfOjZLrqmOzErQZ6JyM8xT9gM3fw86ypYnPBFstPbh2xc79sqWkZ2bybHe7Cq
pPU05RpKDwZJ5Gc84cXKpZPTjMHdwpp+riwTDaMTMPC5HWy3rPiAO9K6bIo/uW6stV47gw2z+RoR
mgy5vv80/zELRAFtnGV3QsqC13QCAWmjRLgFEzAPL8jSnIMdabuFjX2gngqj+qUoe/KXgWN97IiT
lgs7aqqa6sYm2ofiGdCaoMo906HZsE7O4xhvcDUmbcHIuibVPgwOLFjsDpwavvPHLvY0bKrRg1JN
O40GR1Z1RP94+nN9JUqlVo1cJI/j+AK6AK04HKMI+RVVT0Ix6NfjUP3Iw/+MqwzTYiTOGHas0zve
ohLV2mn2lx1uHLCiMhKEBjokjo88NGbECmMBfjDs2nElnNs7BuqZ1F3z2T7k7Amg4M/KHQTkrkGF
NhDhVQgZ8zuOf+C0fWDYEOtMbqHWXlArKl9Bi3v5gS7YNca8WH1RNPnfe7N4TY4VhXtpPTbw8OGa
vs39k6yQ6dsRWnvQCogjdb3jquwlXaEg0kcP9cgxZLCIB0s5lnsp3oHuFNFBNiqbOSzvY9zByelL
VvYDTdHK0V/0TeRk+sSVSg3YJ93OdE3w/+bhTjmjJpPXtHEONTfdxgwo/8ys7etSNlTWH0GeMFcC
1a2pX7GLEFR9Mumiyt+XqjRKYBUTqRcs9OHHQPmCiFwudTjAGAVSi5PJXTz2giWWbPAaB9QwqVwF
ezYiQLi3aQphI0q6dOFcltvAGrAOgvQ3yEfyQ0VFtN36/L3PBYP/UmJACk0upDX2OZravNutEH01
emXgqkefDP1QOYxlwmPL3zFqK0HiKOxNGxXAsVnp+96NVnCXokDOqE9pFaLQcFZFo/cUjQ5XV1b3
fKhMgXlVUIsF+vQ0Re0K8ydLhm3ShjL3G7uiU5T9VbuZdycUKAkV9lZJjM0HCSAQ1RIvn/Cc8kWk
tHaJ/0R2wu6SAPO6piDmqcT1mn/rQVJfGJAO8aCgQHzZCJZW/d31wsaG2w0z6Rlk7e0w1DmyPHTl
ojUkpemTf4SHek5PUpg2xf77DB8HvrdLWVgd2tkYPQndv6oLmEXDqu052iT5oQjHT2BmVkx5xNb9
93s8PLVwIauwDmARLYPt7Y6oqJNKHXm1aVXWDbM1tXI9R6TTqJwa6lcAeFMetgRILRHa1kHJ0+Y3
hqAo8rJBc8dy24M0wKQC6DcSSfsMbNhW49R0q/j0DTzIszL4ygn/KUbbQ5g62u2dGsBSf1FnJ2Ne
CLJC1sCQwAqyZjLbIiorNiw7ypM9sXbhYRBnybEEzGKFNdnIdO2K40TBcwZtxBmhgOj3v214Pb6g
uYLTWnCpHVeghd4+mUpqCotqutX29YE7QkWSlVq3Z6nZgS8DpfdOJwYq1Bad35ZsFQARPE/EFpku
//7lN8N/NHn+MnTMOYC+ZuhLRqQN9A7ipOsXDhh5NXXLSlTB4PGtmfxLLgCVHjGNKZu+z8788gFl
8IqVzKomXonwTDwqvWSzQfmgpcGzx6KlPkoNHp//VwUHHJfha+JeW2mYv/yNHv7CcDD/KU3aO+DQ
rFEYdhgBU3Zeadi/r2F4PxuRlXU4riIGYhcOOuBeB68wBRYle2Kd5B+3HVYsEAsiQzuStuiwQ0jv
lbo0tqLSNiaZolTqKo+0aTd8vv4Cti7A8KSbAqKQfq+phw7FeemLyXkrH4PdXr+lP6zALdJ+89bG
cgSwyPtL7UIcOj1LcOFwgozqVFIuU8VX+Z8pYH/elMTJGciQtlBpUMZKcHq7IejFIHQMK8IjF1zS
NpKZzKFRLwd0cdDPMw9tFvy/awDUkRv5mb3o907J225gsGsBXLh84pnjpMrlxdje3bu/NmFYov9u
zgtf24EIpTsk5FdlhGevn6DTxbRS4Ppmw2hzZaulilmW2mdh36bZws9P/3Tx/lp7YadXK84vjWbO
YB3KR/GlMBYm5BCrWnrYw9jSjTfvLP4rcYL0/qL/Q+OlIdejyBsZ0GITEGOJBvok4UXSnd1mcaos
0+i6lZQm0rOHFW9YTms5d71rF5Yt8m5DN7D33s1R+RP8MtrbmUswqO2CcHzyMEyqHgFcKo+/Xwfl
EowZl0tjLGtfIpKv/gHOeTwdZm7ag+6alWnAXZWjvCVAmh0sf90+1jpHC/lJhCojrBE/xpHilbsK
iMCmpMJCuxPk0e6+Fh5gSTeLRA2ZFeStoMFy+nYiZz3STkDF6tloFdAZyH4FU1UrKw==
`protect end_protected
