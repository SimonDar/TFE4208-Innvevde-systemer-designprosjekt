-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
B0GBwSbvMUx8mH5106Qe8yCRdeyZSrorg3UXbikBlqRiWjHGacl92WzC6TyG24Gn4IFR3bRtOoY4
fAPgGBirlxcygWu5sEPhoAU65gcIPyJaLPya09RLCWnHlfY81fO8nY5kgy3A+gKP5CQdm4fg7daA
ng9EC2CnCpYXEF6hGg3rZXzXGPCfrz3YdLMn/0G+KBdwzOvd4fwmN247Y0pToHfFkXC/I2eMJeyt
KdWLXv/5dM8pnRvScsx+plJTr3bQ9OxgnMppF5KNYJA+qfgFU8TzTIx3kThqgUVbAz1DVnJh3s+K
SuvTj9Hf/MERTxbxlb1TJZwXvLDV52nPluLk8A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
Uy/kfyYgODHukVI+6ZYGV6g93H2cWXrzZAi9jKeHNkUeP6Y3R7XkzFEjxjf01WdU70uAZnUgqT6B
J0Hdzwm/2cnis9lI3UAP3SolvBwzPWVFcVa8Ovit0VerJaNuaHpeXVi19itGS4lAJRRezYCA70Mu
vXBIqrYB4Zf6IfgnlntZH3YiIG48fApb5C6Fl4FNdhqweGdunWCJ2HbJ50Ck69cdKES08oj0LM0I
0cq2VKyM0dYBZm+sKB419WI8kbnOB+XTY3XWurEL1BcVKZxOQSV59g5Jz6nt/PmY+aMEnq5MTWSn
qj4M00Fp3P+3Eg4iIXBBlwXOpTOPkanuIaDnP8X59xS+Y5IHLDj469o2XGqc0G+am0QIiNKfKPgO
SgT4SVtlcxf7F5VM9DUMEL8l7otufxf2QMI9iQdWkPpwzO5ywoiO2gV8a5QJh03YdesBb67ECO5M
uLQ8zuL2J8bK/zdKB9nD9NRkzPilFLr5KdCQG/3J8fHcqYdy95o7rgyfJHgETiQeEOI9neDjkttK
+Gj6NgnBkj+4+lJuqr2Bz82fFLZV8lw4J1+URiSEpKUOSMvL0cTBqV7IcB37cbHFIdX3twZh+rC6
SMPNRHyLmtiN3750eob1gdeKVI3DxcOlr+B1ewalotJQdpZqIj2Z6UX8of7lPpfVT601HQSwc9r2
y1t1NfIbosf/3z7HUDqsmyVAsxGrwIGkMupXmi/WawxVw/8YWrgTcg8hqq/bMRO9jerUxvDAheK6
+m/EEWPcsB53xAUD7+g5BkUorK7XExBcmPU09nGrmp33a0kRV5rtBBJJlMQULUWMnPqHZ2AgJmJb
SX7XWvMNdlww+O4H1+UzvWVFfxDtJu6/XjMe+cAL6LBv2A8XxXeTuFvH2ETh9cNt9BwQgU6m8vaI
V77gou90LlNCSAq8PnUTjXGvQBq8UmDARhcBWPqkCAWY6I1kYUn0u5L8Q7+XoDsy5DnWZNFJIXFu
R5BTJVqi4SRX0bmIhMp/i+ipcojuA63eciGqixOfCKFromt9WzIzv8q5OQv0ZuDfdnAvYRuOZSOn
FKR/efjaNgbN23us4Tvk/Yv8wEDIl4F71stZP6/qnZd79+F/tO+kYHI2f0hJRP5Af/mVIiOanwEX
gVM4AJtQZc4ZX69xbg7jwK1ZNz8PG3nfHdDsTkqrnANEUGTE4IUQgw4bG0NRxA6OZ84yfEGQMpQW
kTaoPj4sZBaNpKvdQiNR10unFAIiR+c0rj+VwN3DMPAfVdb5FDkKOA1pnNWy7pcjHCpSJDN2w8AU
M3k2yuqnGXRkjZ127dU3XSbbLyaav6pRB+SaSX7Ydm9m0QgfU/lad6904UEsse47Ie3V7BH98Lcf
zd9Hcv7nKoKJttcrMxMfogbo2JwCjtpgacT9d2qTLnpukQE4e+9qRKcmrya2ylSVqULxI0fALyec
haGsLR9AktBx1s2WpDQIE49c7q5b+r4XgM6ru03RUp9rdaMDWizTqx+Q/gQ6IgxjpeTvp4sBnKwj
6Ws/L+jmI8YuyPZBsYtkrY7oI/oopb1niS6f5xKLbgNnlcZ1Bs8/tmmuI2je/W2ayu7eRgnWIQkw
14sXKS/aZJQQn12ehBXYKMUlQba1g3QbL+zA3Fbpm1nJmi+uJiNVUIIso+U7sv8DksIDcWasiA1D
gGuU/6W2j+jruSjchWB/pON3ZhtotcxMSw9hSoxHwJPuU4UooUWzFhPT6yEWNW+fxkf+dhMXUUWC
qh9cMZUt5F+6g5LRL5s9F3tx19hcfaXphoe61zwNdavQ7WUCUGOZpTwPEWkBEGZKzbayoazsqp6N
07MrUZ+zCVsSN3owYcr0hgUuhGJYcJRc4zYIuo688P9NkEghoR77opKYfcrINMahwQLDCOIWcWor
408z/uiCSsfD2nuyPRdSl8s3i6UiNZQHemxnF6jlGPW0JVcPB7f9EFJwQEuOv0oh7KLDhjHFytgA
4oCSei8FNpQaGrW/4xLtBXJPh3jwQLZSzhIQUf/ZQnCSl0eQgciBohiFRCT/oj+KHKp005RX5TlK
mbJA6KZ9TEm0pg1G/Rc2Gh4lSKfijEvjaXxDzOdQPB1hICXHnsAWpaSb8Q3VMLh9Aqrv8eWdHHEq
jfnQXRs8hsFmmfeR44wIMPfVSH4kpMojoOPkJGRNFJaBJQ6DMRhz3eVhmeBFdpGOLC2/ZmlFkYZv
O8FYpzbUX1rMK6DL9cfmvnEN7jb5MuBEzwGfwM+ltGv+chJfZ7S2VLEONzV92jDF7f8CA8IhmIb8
bA2+jJBDjlteNPOwUmrwB69lbrBjkGKm0vPoyX+ASHlHd3Y8QxbUqYna+HHXXxSwEleJ+7hQ6ELd
cUP0m21g7CMWSscoqOxT7cJjpFFD46fOj7EZd8sTDiyYMapziyCmEDj+olcpG15nDE2tJ+nYnn+b
b2gT5U+taEfmGtYoSVQ3eDItlUviWVwpIIgYV9DidbLwfeXKo4We+dZDkZ21n12kAKShXe03YFvH
DxcPZRtNpRNh67qopyeqOwfJeP2mIK2ji6Vr+nxysY11veWfHJ5mF07WEcnCYEQTkE0EY2uIaUuo
8efE68VBYDYbJsKNdDhd/71hj+20fniV10hI22hhYVEVAN4k1sdPbKvmt/Fwf4BCMaZ0bfhdgwAX
j7ZSuF2WHsPxAqDRVPp1390BLZWamk0Ts5wTfVfSRTh7Q5Lszikx54GGNlGjqmdAFz5x2FyMMTEE
ec6ADbzVAXjJibMS7vjF6yRmHExStl7g9R/kKuW14ZLLfLLJkWroABTP840NX0GtueNU8i6xwH0u
5poI//mQlnCcWAg8iGA4S9n5gFlC4BII/g2Hwov7GlGmtGw9t5SYaF5i/nPeLgFXKQvxU18ITP5V
Kxon98jEUM6G33yknw84vWbQdYUjGm9IpUgpnvms617tOunP0nxZTtN3VCklYwIIlDg2cJaKugjt
m9fds/bl+e1kggRTvmOEjpCDZM7a84iv6gJweg2Fhsf5uCPjazmPY/f11GriIK9NfXp8Lby40dhr
AuqmhhmNHOFPUy6sxszBTScqGUCuvqCu4KkzBWZQC0Qq1dLscRs2bP+hyu3De5SyKfpiIgtSaJtw
eql7Ev/XyDK62cqyRocgHvOtzNIJ+D/D73u5OLNY6JDKNQdE0DnwKGrTO3kKaFFVoeKscaotTVG/
xbCZTm+z5sM4PtdOzE17FdJyrPBRvpKA7FDholO8fPcgczhqoQk+SQwDy2Og9hCanagO7q74MIpd
fFMopM/Shppvy8EJgta/s+CCfyd2NoQiZF8BuTSbT9z+47z7ORRtobdK7vEi9hSbup1tKpQ+JD6Y
lTchiD8Lfmwque674SV6dfYdnA2dOgdcZUQXJqHjM/ef//yEK1poq7vL7DxHeEGUEB9y+qV8qRfj
yhqv90d2nqoTiF/PdaH5CWv+UeU+yFHzzyhTSHTWRQV1kQtWCdhjKHid5hSMy3p9lPhm5BAUHn7C
LOva996PKT4NBzO5hoXTSVR2RzZPo+wYABEpCv6a7axu+EyRTrTzH2bgaqbMKp44Uvd9vXnbH5wL
XvITkYeWDtg1z/ipunvbq7CTIYZjpGwYogr+0FqZ9m6ZrS+C6kYCiwO8JeSOu6uZWuEQ42n/tjay
gfRAguNh/Sbh2CaFJXuvvSaQ8wymUFGdldBwD817nDlM3Me2xtGsFVYM/RPTmqCn0bHKt/cVtpD2
W12h9tjgb4B72AbeqzyUmTDWrguS5XBlarvGkdYULMIDp54wQ/vnoMHsewZfridbPZm2c7sBAh7F
wfTQ0cxtPquDEdwycnM4q7rmC7B9QUuhLQYsy/rHzyVsN37lbt0ZqJNrdbw1Q04TiMoyQVVuPUh4
Nkf6YzUdsb2+iyxM+Qhz5CFzlQrfqy53U2Qhi4602nxrNb5poREUUm3od3jS2pRzn5KQGakargjJ
ZliNbBojyao5ss3FvWH9Qei7GaoxOPYsHd9c8SxAdsLRDDKRisiMvwroLxJBdrpHisYTXJLxcnqt
Hpd1H2wJSADfhrtnu2kIAuzNrKbkcmPCcxDYe6O8n7llRFFBQiCRm4Y1GCbRDX5rl6L9mgt+UP2b
Rwsf7JdRZ25pb/PbTSRXKFBUN0dBlUCmGWjP/ssHkRM/1QfvxNJQPm4hiL+uMemgKg1LkmRWgu0A
QvhozWF0fgMZF+i2fgq+VJToZql8K34Nlvixi91dZiUDgpkWlSwsM2prMYWMcVSJ1QOdP7GGVeHK
EyDvQgBx6Fon3EzahXy9xNAO8D+r7/aRXZ5c49di1CBTBcu963Pxir0RQVREZINOCls6GVabmAmh
oDRJao9jWCA4s45fOUDtKB3kkErvipHYJfkVcebnHNTsB5K5YnhSG4PZQr8yrbNAeaVJ3bzWF7yv
t07Twb0/VfBvZICUHVxD7QL0SCycXRT2csFlL15pi4Mq3nFEY6qjWYuvuzidoGU2GV2dFvh2dcoK
khIIEQu5ZBzLSnHIb7QF/tY3V49JBSI2CEtLfQGMKMLZd9e0OYR027bmtd0/dL5NdzW4qUpoXGKY
SyOsXkaSkGOKQpBV6te2/0IKOaifUMMC+kxFmNmVZil0v2ffDHTnDbAJ/0/Bvcqsh241b+n5bijA
ZZzmuyDpKQSOshb8oZ6A8M4tmErNdYVk7abuLlnaUPB99MqrelprzSTGnsDu7Wpf/V9A9haEvhUR
Sn2+4GMUgxm7zF53/O/Rkno59x5QmkNcyLPvZPUfSzvngmBvUt1KUvdDl+avLwDIxpROAfHrrQW/
E3y9C0IjMi4Xk9Pku1wrEWQxsbgSrUzDKR+P8kEpXFGPAumyAYM5RJpn9dcYwfQTYC209rIdxgNA
aZwJcAQELx2uLVeqP0utKdp9Jts83VgeWNwxTyr1er2Vwwp0Z5pHeK37SgfSoM0pDRJiM6LwmhTQ
0+s9VF+rlBO6/g+BwsnC0yf7HKdFIky1FAPs3LQwZQUrc5QTU/QDjlj1FzNS3Jjz5FSdVHaW6YnP
cbBGc/Zsb9F0Z3I4XZD29dIwaHfLS6Ow+MON+bbN+YvtTqFVYUdaheK6Sauem4f2blUY/y+Tg/Y5
TWCBIZNmLVJMdgLck2DzWbL6IbVjZ4hYGGZFk+KXMcsOU04Uayak+M7Mf99rfmSNU7V0+HRH9BBh
UeHvPW6oudKl4L523H1i2Jz/mG3l8Nvred47l29sFH3XLjSXacLlPb8dpifnTkV+pIrKAkGNq4VI
EYBk2G+0QBVtlYJLGkcPnE7BqckPFK4pnWFVb/EZURCj9ykvSbbGDywrp/vmfNmotr0YmwMvQorn
z9uWN+bem4yNQYND4zTzjLvzbtIvtAkwdOPEfVn5vEmQbufNvnwAvN2T0hjRmra0PQ8mTjj9aq07
uWfaJgXrrnJxhQ/TwcBFx9U70/Clc6YIMSFBhPpc0SnRCPyxYEzQ2Rntasw+yHLQE6cSEnpvdP37
M4k97n9ZCQc0g08KAz7rP+nAx3QNYE5GluUxZ8bFlIR0SfWB4r4wthpnyluMIdNNtMZRDt1iDuYr
X7WVOzVyCjpeBQh9w/3lE5+Eon+xFwWd7BKRLWI3HphpnQpB9YjKwgcR4O1Uf+d59K6/lXOBXrc4
3porTVkwuc0A1NQ5mM8gD43d8oKEX0sQ1FeMSm7miXegGvkym9Jn7pmqPj+hKSWwiYMGgS0yRWYL
6H6oDBgVml9R9XVP7L1rr/W19UL7zz1oWyTxVjaky2/qPzxYez5t4s3ob5bg8N6VjpunsTLVRU87
0PaK6d60OdhoGcg/Ah3EduguNjfjNEqKimNl0nGrGOwjHpfZ1+yClNbfVsSE0PDP0skGgJABs/2/
65mzVmCyBa6Bk75avuC9VjSUNhXKD7Ww0RKERjI/gWRH3uY/6BMRfTKSx/Z7nTzffF/V3KZWgjPF
GNLh85f4EAjHLeUaX37joVADDQg5aRCGvETcYhTIdE2r1sL2K+dv3JrNzvtffaUpJNFWNwFWvL4g
l7vGJ/p7qM2uEbuPFkkd1PPsCxbWZUX/nQjrv3Tu5kiHRvxtSGxVve67UHHtMAWvdOD354JPNyuh
p/tUHcSgJDhYJGF5bC0BuDz5Sa0PumLZgWfv6AFSnUbfGySqTTwFeIJLKFKkz1fQQA1N6OXJyVQe
N+2N5xpMUgcEaYHQQFFBrt3uVBFwasXnaSQrzBE0FaieGU6C2tlnVR9cwoIFLPaKoaZ2LgLNkTsv
M31iGx7y8rx16+I1rSC7rWJK3F8pZh39LqIX8nmnS20vszeKkR5NU02dmC16cNO8aqQm05OfteI1
QnDxSqBnyHKms71e/94GqdacZVzNH/jXQG6P+Ly5B1zWXgAy+2n5fJA6Y2ZNGhYuAQqmVuBxKoIa
VWDZF2h4La02JM68KiUsefySBz5SevrksSQMroayR2hrGUqRBjOP/LvzuD1hOZz5sGp+HM+cmUqP
SZnBaD4fYc8chUgjzk0bOYdPByD/SaQLZcvrk1rn1CwLiSc9KVSfVs8N1FccVm0/G2NN1LJBdKz7
4bWwbvZVp0Ky7FtkG1JZVmoIE72AgJ7bPfcW3VW+GsTrvHylMeVvMY4ELsnpEyIEImf8s5L7uJu/
vzIs3kDYveL4R8QcbNmfnOdt0Y3Yy8sPsZ1rDEX7OZZGOYnb0sJn7PV1HGrkobRzf0Lwuw6Zx5Kb
XPNzgBOYi1fggCShb5eqbPs7ZN8SS2d3i89DxThYT2+biaUUfiXB5oxcLYYKZetg/mT0q58+H52Q
8nSucxjrphLnpvvrhuzP1M2FJTn9P/QaE0yBeR/aP0i4pN6YvtU4ro22+0+pI1KlYmcC0aF0C6g0
LT3GVvIEepAl4zwiOuHoyUTTU8IGYl4gIotLVIyJCtLRu0NNtTQZoyiRLc0ALCBknbOMk6NwEm63
rc+OPPxWbmljDphmwdSsxyxxEYjSmwBliIzMIbZ7C4hpSbvenIHSpN5KWAepr193ucAFBY2LbVlU
1FgYAlqmRgc/2vWzUMvU4+xL75MXDtJuqMG1aIKiZG157ilsKE9Ql7V3x7QIfKW5oPZdRf2fuZ4G
pypKVMdeaDg6avs/KjfiYEK8BJb9sqMBX6r3FOUvH7Czrx0bNDCQ7wXOQZxtmbc8a0Y7BTbvRhTa
KZCrr9x9x4IQjAW6ZTFhX6lsjOtxmFWZwbmCs5my2diPJHySNKWr+r0XXXr8fC2LJ7YLpUBzPd7V
ir+rgHj/pQviZq/wOD+eB4TZmzVmhhqBmy9QSAUSWwXT0iaQnjIqN+RA8sA7WKqJc3Gktu1BwpqG
owhPUuMQYERuvG2vPg9A4NXaB2UyJMHiDrQBIWfT59/TqYXcqlnrUrMhJMa9Da2UzegM7PKocEP3
0J2mjFQ/w/xF6F1rwW2blxQRPa+MwW5jGVs19eY7B30gKlwBvA++oKnZi70q8Q6E1RTPMjd8ojlW
fvpAYx2tMo9astHAy23+ShlbuoSoHq0jajRMbxLYEwEFqErSjxX0xc+IfhH2S/g1xyCRggZ/XjQs
o4b/F79Hb9YNYu7qGioAbdQaOTEptiwINCzt+VYnixWTibZwvQugHtRBrwaj765jvhh8giTpUuy3
sGN3vcyRHBIaqLIU8HX6le9lBOv+QH8Z7A1D61Zh4mg69SQpYuGd7cVYnZqDoZTZ8Fc4jMxFf4j1
5M9rr8Mz5m9q9bhIEffGLoJMWAr/qWtS95ZWgzHfIJSS+meKvt4dWG0V1ES+j8Bb8su/R+b7QkuV
WtodQt3H/62NA6rAeFKAZjhT+2wC2ZCjPvTOCTkKZ1lGiG5j2NhCeG+ENDMsQKsEjWoEg/n0CsSU
wsk+Ggo+H3sd3+8UcHyhodfkaB0qEfZy2mAEXKvliVJCAhHY6sGP8Vf+eSXNpbOdBM0Gds/yzHkw
SkkQPnZnath9XXHZFuSWFJSe+7adnG3XYL2l4mBLrWBIw4UnAbHBEyqiM9Qn8QsO7NVBkfwuFv7D
H8MmEStXisD0g530BiPZNmM85nqNw80+SZH3+38VfjdL/eVaAIUt71qK3NYk3BBkmd3BAH7h+jd1
S1qmR+hMcxjwj9vlDKBN5obA7VPZOwUg9MEDceJtVe6Qg6EWNrourGhtB3gtqLJIUUSa6ay7mVCl
h01pNasz/gS9Qbj+hZvLOkdIzppd37cuoUHKdPA2uARdkDQHeYSGC9LZbtRU9sIT3Td38iSpFAIf
UyQMP00LCj8YP6xMrbJfbMS+ECv1XQXvuRznkI30ksQk/lrxuTkRsbKmagOblERj3pTAelXTvLIp
PAKtGDzVaLV7n2jSBk2zwlP5r4cLozrDBKqKltGPR9SuzF/B+liLH/cskWJEUTy558/lVBcW1mUr
/qAY4RHZEUUB/5f4TsNSSjJyiRF8Oye4fDfLQIRTPGXzwQrukK60M/rcnRp5QvYsAJjZu0ib7IPy
wLKGj6cwRU2fokVbnmGHFJu91oYt/VG+8qf+ePTt41WlBuGPlVEVX31KNruo2WLLEim7NXGPVCUB
8tiAgC0kNx0LJvFIA5fpp0dwaXP7zAQc7qdgPTSFq9HVgkbfoWtMQuYgJLWX7u6QpErB3TtqyaC2
j4u1zUbmwVTtwYiuperMClx4Q3/tUMw/VzbMbiRUMHYlXYOhYfI6qCA14JVsVmdiGfAlVzmEjm8R
dKaHVCtxOEzH4lTTohdnFrtZP1MDUHI6ZsswFW300/q7B6FfRnmGf4Id85aZpn977qVes+fD7nu0
AIG1hX/LCs9tboLCh2Jh4THt8i0stkrEhrcAU8IKTMJxzAiUnk3wxA71jMAtLOVbhhIiRmdaDYC7
yzHWcD5JURu/lk/eu1dtHeQOsAzesewX0AGjsrnh1asVnQbvYepGVTVKXQdiqKGvjpkhT3Uzlm5F
okjLKXCTZgNmWLacz7Ii2S28vcXaLAmNGpufgAfUlAXqFGGDZcSbrifMnh4Pwm0klsoi8305pCBn
io6jl0aA6VSXXxZ8FuW3Xw/zFKVb61SRuqzux7z0Z3SCdCZz3w0V6LGy7rTbrFU5QOjoHXp9mJhq
1bx+QYRLP7lLFjeZ17Pf/fE9n8ol4N4CfURr+lNvqS8QX1yTVAMjppUGntQlzpet4kUvGpHKQ95F
TAgL80D130KTGL9WIL9E4jM4voy8fb/PRt94M2BiBbL5RDAH5B/Ba8+PE5qEwsRvWqSvYNu132lG
ZgtPoNdnOEgxNl7KzrO8aibUpShk9udoDDGWjpVBwhomcn3RJ3OyQTXmoaI0wAXqmSDy5Qqr5uxr
rS/6LOyO4g4cHjMGXRAsXWPmCA1cJA8+8dhpaqBOOqTqc6T0lVvMz1v0C5lxofDR2dN9fsyGvjii
5AQJt7yqdSs6rs5cLiXtx3XXBnJFGrniZBeqSqo5Ym5Ut+uNOsFzFYrVUktFc0L6fKDWS3YVpz/3
ZTK3H/MfYQrEdafgyAriAXjomxTsXEZBRMhGmRITRjuQr9WVM2xri5MlwDVhLTMrNP0STZWJZG4U
uIsoCihVth9i1t2nKq9Vp4EwHFVwCStH7cORMQ8dKg4rE99Xw9wJHmmNLofoTZ5xiXMSgyfiOhbj
xcqZIpfqPi0mqcjykfnfeb1Xbfl0IaR/hruMJUTTI0Lxy+D6UCgTtc5lVhO1kEpNH7WGFsOM+hlz
mnabrBeBZA8CUz0Y4GxO316x5g9VNADhYNGfGP8BeySImTI7OjOacxir0NbdePwqgXxeI4quXRS9
ybqnijdIDcycCqpcnarqXihX2mRwISrYM/V04sh9ju5OL7tn1zck8eBH00w1PCn4HhRTyY+zV51E
66zKphh1Squ5g6obFWytpmVu623xNdysNrFZce0ivuFbNbZhEWQ81OGYudEEA+gryg6DYBzN4Vkn
uLw02YetWt9U5Z9MaRNBccuvUEhDwwF8O08hIJiv6uEWPc025tkPiazunWu3P2VxDe15Cu3/tGwY
ZPrn71ZWbY0LNy7n1Vh21KIbbd0jSbSScTC/e+0MEKkHaek0HtONN+WWgnWhGn0raXIVtw+JmOaI
rws4Pvsb/bW77ksxvQiQwkVomKL74cE84z3ES9S1hcmkRCO0/etyqC0G5VxtaC1FBxSRai3SVBEq
U2U+f1XwTiGxF8hweJVQPRKIS4qtAZrORwC8c66RuAL1bEJwK3/VnycY+uMQs8UrvczoNxdAW37x
ytNhhjIf9IGwv66csbdQk6dwgateOrIEJ+TfXYGmpY3erpeyW1pmR0U7D7OIRLjFNn4YFYz7n5F8
McH2f+Tz357uHmgrPzINokbERdn8sD9nrBEm682SwVBOWlH0OD2rfDEFXAKKUs4c8Z9Dq3k5GDi4
kluLGUcn2v2sTfWFIygrHchBRD8nVvKmTAgYEB62PFSX6c3DZFKblDfWTulLrxVclrCSKcNC++6j
k1u03vULa1m/OtC4PUWVYQqOLPEZgu77rcygTtph1hfnB4EOsQpaRXHgA0KjRAYfHcXwRHwxkjJb
cJs1D98yCL/jFITkugLdBRHT64l3A42VLPMijGVhx+9Sveo4vcbW6gAgasw3wtOFwWS6gYAhe183
oS69XN9EgtkcSmZlvhSPcYix+UP7/xIsgrecn8avqskUuiLO4aTCQJme78aIJVJMpwATm2Nwkgmn
DjOP/sxoDBesDDcaqVXgBcQbU6nH3fpljCqOT2YxsibIlZ+Cb4YF8PSdL5wPeODHI2Av9hJWDeDA
xUmzVNVTWURahrhSIeGAOalsOLxrpO5FS8c7ICQDdnCZlaIKxluKt6PpufHID0MuWhUxmzxxjx7a
6bWSuXfQIVHalIwHEBoXp03Tt3H53r/BvdVX0QQ75lInTA/O8UPNmdHKpq71V4Li5q3ln215psuo
ghsv8Yjby149rWzcSmwc5abkwM3hMh+U2IbbASM+ODCzGhn5vITE28HE8c4Rh/XlOTqys/vuAPDO
7Rz/EPGU1cM3zydZFJNOcRqKDjnACDZm+heaOL9GgCoC+bNLzV+e5GL/oD+Aj3XBF+tSEF7A67w1
VSZf+0Lx8uAOsLXr837Mej4Z0HtRnAHzqQVOb2/dX3iGF2j2HrbEyQY/4qMbILaxulKHUsMwX3nK
rDsBxHKFRfo/9AWSYmV4YUaByWE3CdZBZdZkNleVRLo60xR0G6ZwfiIr4zwhasJ65FrPDeA8qZKw
AyLrbx0jNet3AQTUIH9tZfg2Bt+EkLLz/a2exRptwdmsUPBEZFzIl3kINLCz9dC2zhiJrxBILcfB
NEhz3BE8MpZAqN48dcs0ZbaF1hL5Dz7S5t33lXPokFDe63tc81bMV50u0R3ZB3bfmlevTV+W8OZf
S5YKa+ExLNiWU3k7dEkySY4guYNYx3ml2zWSZIBzjxhK5OFJuRLCWOc4URda7v4sv2+XvXFA/jVL
EfJcNJFRIEkQt+B/3sa0+NSGjyfvl2MzeAYgJuFkbOEdnO+FwrfNP+LFtlA8C0graVihnJvuvkS9
iq5XUDHA+sMw3/8SFFVTJS1dsjiyCXIdLUQO73dlawKzztmyWSCB/yMIcPbNhBIiqPb9fTSEF6xD
ybzzOkke8EBWPLq8WO4PDay6TapmNpEie1mmbb4W43kaFj06lRNOuBKXMj0jtjqwwgwW2qQf7cel
rjmSXDKwunIydz5fXHiWgoWCNdgaPjiBjadkSzhTMUArovm6zQqHSO5GmK7irLt10nuV0J3B/szR
bNj+1zxAMPtxuuLmHiny1IQdPqU1qlimD/g/n0F6iTqTqBwbBctuUrzNRqkLLEnL6+t41+2yXK5J
C0m9CEvIo0IO76MafYjRjS0MQ4sxsnNuYW6JRUKQLPXjh4U0y/xSQBBJJCKfdQLziY+i+kP/Rvsf
Fc2wYSYzQ8sqMpx0VSwZzuar1PiipwpKBzZuemv/ghmjjgPJh6THUeZgoAsRFWVQ6BU7A246x0Xa
eh6hslCQmb2xDxPXQXjN+R7qAhOt7JvrbtMq7R1FXB1kvTxhPhkTjkxI/y69CQdXNeBSaXHvgTB7
uqIwBgryJfqD+6iX/z37DslEXEK3pjDUlo/6Itt3J/Sbt680eKOr8yawnogPpfVlZlrdWAjqsUKZ
rv2+9a7/KDNt+lF3s+ehykUM6CjHpa2Arz/TcIeiGaA+ig9NH7614ELM1ODAR9dDTCOUDATCAiFo
am9NXJW/n4hvK5Er4b3RaJ7pUADUmeO2in71FTlEqnuusXDJtbHaquAHqUzsdeeXgtpUWpRfMZjR
SS86lNrB2tjxk1d5v7dm60lJ7X3GAKqPNkpadRbEGUju/KVOoacgvQYYlRle60tpJjUpDKlZ3ztw
NZvVHgabCR4cotLtkuOEue3yGwkHI3S7lLHNI8D6y2x86E/3wsdIf4n+YcK3nHMYF2xZlGrYp0bX
Q2wK0dhGwc+YCJaqX5ZSVEvDBtVDMQkeCfLhdpt/JE4l4hORJ9FuRxAS1AcdqB6Uopvuyj6zrA5k
a/Hb+4NeCuiW+LSmh847N9+DJUhmVzZDe0SdZXMb/Q2myKXKd3/1VgZn6i5UIErOCB4All85/sIV
LoV3WFtwog+G8OYdVReQVPVstB106zfvkbHN7ZjUDttQmn/phphJeGlN2sRM5ib7op/pxjPnWZ0u
ukYKxyFhcqtWQ+oD4rVEkN+ewYv17vShtwuWILc+uaHa4sZxTBqF2XgOfe53q4PEtI5dCrRy/Nfl
aK0EnSpcaIjRzxFQY7RaxSJnSXsPqoioor1B3C5T56hB1bsyRLgtfIyc9GPutabkK5CJejWdt10y
t/xkVGmZyQPC53Z8vJQMid7CiKYrEeXy5lFhBPxUzRLWfC21coFBkexXqKQOk8eG6pTHSctLpud1
r77Bp5w/QJuLtn1Q1U1BBzF0nVnm+55HqUapvjc7kKzF3gFfm3zfBeow1NlL/u05jCvZtx+2z01O
6SQ0UtIg1HedHwAwcqapEmiCqkB7Hg==
`protect end_protected
