-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QtOmKyq01DRaZSSs68Wjbo4G4597VofvJg29e+fKrfX4VEozEpskf95td20NbYeBf6h04bBwo1Mj
+AWf6N870Iz9AUfbPH0HvGbqVs9fb9RzRNvtiPrABDhJMlkFcV9ulWyx97A4VyxpmT+zJj+41y4l
OJezMQB7bAhnxHd+gtgZwB1j9tq92osHqNNk5J4juvBfKMl8gyhP9vAUdnM3jf233EYJFkCyfbwr
+o6TAIerRkDuzmRGZWg9Mo9kUJZljYn0f8kqNyhVFo/YiPYAbxZnbmQhni0w4U5cvKcWF6PiVQdD
0aZEeA35JqnmYbqblEA8hKFpXJ0HVNRqKlWeQw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
qRGPzvGXd3+trFaNmnfw1Hk+wodRH7XGYyAh0TPdnKT6j9wwkQVxdz3U765IEsxOX5Hr55WwgYZm
pgUNrX4k6Bu/cs1oNQNjvdnjycCDYZrifz6IWHOK/yhBTxvToyFVXi0QouG0S9g0OkgaJyEvY9cn
00k+py/4T2nOkEKF/u9DxCgKs1fpMbZ0lfSSspp9afK8toYERaS3oa6CdHAmrQCEMbH7V2fqyk7x
Q/1lUml3CgVWOl7LrlzJK9UMLm7V38UAlTNGvY9CZ1LPX+UgdDIO2QG1oJ6vbmvANxewQHWgXx06
gVc9eRDHkPeG7/8OA8f8Ia8hyXi1beZAsaiPq8UJm7/azpMFxjUXRgN6DfR60XV/+Uss1kz52pwB
wRd9YJMeuPO/dREt/O4N6PEXZETsuKBgu1QiHQ5FFV0lHAcsrTM51Yzslxyr/TCwc+OvbXKgP/z5
C050dg6qkeklqhaDY/ME4As3aNUE3af4ldWDONZbewhjH76yGvjEWgQ6aZE6F78RqDVPbuwWjPWQ
oD6CXMMaiHSp/rXC+79rE2ZH1FbHX1GcFc8X1OaL1vvxwhkPMP9hJ+aaO9sQt5S/x8Jz9SnFPttc
cHo8SeY52gfhAG9IWl3UsUSAvHD4MulwUYi+Nq5FF+RahPZtma/EbDT1FMH0YF01VdniXCzgaymR
dg6tlZAZSYBqL+T/YLmgkbMqmThah1d6e03U7Et61X+40jOzdBWC5e8t+RQ9T79m8FPJAGcdn/bI
X3AjVsMPqvqzbjyEmeiMOdrsc2LIcmJMwFylX49rwzJYb6LbQqpSYim8ORLW2nkm5YSvalFiRzKR
l6xKfb/cEYobZ+6m3x/UO0xzxbHdvYcs/HJBjfPyLkpnCrU8cPry9nbXWWTd876uXsX30/Q43eqQ
AQOSPsZlr50tq+qsIjvyKNo6TQmVqKM3Ntv5uLquENdg/++O3z+rF6LbH00DOVhincI2oH9obXRq
Z82nC74sQij8bLes5GreVO6N9wP3NATogy+DIuMWb20JcOiHiyvFLRFuBYtsryBZy2+la86cEy8v
4sm8eIk6eI3XXKY13UTi3JS3rLLvV5KBP4LPz3i7B1FyLwZ+0pkQffjuHm+W39QyDY/wok/X7lT9
5k8EfbFnGZ4VvTDGRLvSt7Mt8xp7hkrI71yzHd1p50+v0Avi5+NHryktB0spjqUdMjhodwgbMBTh
sHBQ0xjK9xonpDnbsY9zIEMstahfjjxT4SD3iJdLS++TLHbdGupWFB+owa4MDzfg0+Jt9KbfIL0r
2TVDwap5CmbGgYPwRh22tz0ER2Tv6EAOuDUEwvxCp4Joil074DD3ywbrdebhPeaukZ8L1vtM2vLk
dNi3uxzGuCTyn1J7sQN76ZJ/HpUmDu6fvr5xe2F9zgpJFuX1Qww28wNlGcfMBNZvniVcntbU19ub
VvEiW28ILkAaEIA4zwn3VeiTqDJdVsvj+FqLYT1/N4qpaT6WaHvtlnREUY4TB4naXtBH4whc0GgN
7+O3TdYLdSgk7cLidkXi1Hh3/2me1zc+uiBv66CZ05lPPav+cc0MEtRiAScYFnzW3fs0G8O4FUX6
vdLchWGOB+hg8RAxbVySKlUL77AhT2nJeMo4UOiJlkX1nnFKaGeZC2wVvHRRg0qPQ+XsgxGAb4XW
2/K8Ad/rx5ejtVniQedyT+UU8WaAoSr17s9n25HZF3zw6jp/W1cXrnprSB/I/DCAczhR5577xfT5
KRAIwVGGXkoZ4HJTjGy56e7srfjdkNWyTrgfPnrQBYoIyDDD4x8596VQMmNTgPETMKINZWKqHclh
0AhJ1+yJgxwJOqUW8czU0MGpy5S7xmG5kqYMzeAlYy0tXWEyaCeEGO1wdfZwlMzaT73nP20BObEI
YlPAztX/Y5cfFAx5cog/gwN+uhuH2g2hPujufhc7NxQjvKzcTArklyXpAnVV9fz3xMF8dahC8F7R
C/fBIO5dFgQ+EcOJvRvZFN6DeZPH48Qj5aYrQwvsHYHdILhO7hH56Oth/7idgEazl41n2QGqmQuf
2ZKA2QsXmQOor2SWH0a9cn/p688qF6LJ21Bgax3ARBgHtu1ez17auxA6XtIT+9mzTJo2JSl0BArL
yTI4bfHtKCvrtzvsoeGB9K4LaaHE9K7eDREtxG3VY25tkvza2gcPgjMLg3z1xLhhLQKcdxShVk1R
sSix6wJsJDK5ErhFbHZpJ33Nx3RuW8cKNbjtHRhlNFfWWrmCP6LeHJQEg+mKaxi7GcTMbN65OK+Q
N/r1VdXBOs0FEOYILqMfXCFkQd3jDts15DYO+wimR41BPeU1M5NPO4kFKe6Oc/FBYDlGugwN3l07
uAlq6QbduL5nj8KA8hbkzzE3DN+cE+W+otiNlRMWlWyS1zNPxHh6NY9hepvrMxOOewZgTJDdsEeA
XVI17ApfwdvJBHpqlApSB5nt9QLNbWjrj004QZNCWoZEXdFVuXYSRd2v0qo7t2+KkBC27IV/YyIN
cvR/+FK7k4VOZOnEfyBuCd7NskLl7imWY3Df1BRS5QZrsD68cyFEiWXr9hviNOULX9nTZRLJjhtc
TBX/bFXHp+G17EDh27qyXXJoKaX3W/lZQW2UAkLSVDcdC2ou9yNqgw1Jn2TQ6Ai+vo9pv6O+6W1r
Q+68YuRMHKFfS+5941m/4fq2288KWbITRBgrf3KQYBqmtBTQQYQYIeP2HoT0yJOEd2/QuFAfdhRw
QOpCQ6G7c+9zYa0YNTONu+6UCoT045L7TY5T/uz6ptkGvae+j5G96IU2zfMS7QckVicnwtKKtvZl
/keKux5ekB9Y1TGTXOHTfM5ZmwWNEd/wN0xx/U75xk50ZNRv+gzq+NH1V0BaoBWMH4IQapfGQa/J
6M9K1vooMZ3VjZVmMczIG0E7YaT36cGzmz7FpcL0xslIW2nAw3Ig332RSuZb9tVzdxI8O30Bt78U
N8SfEpShffhr37R4+UB6Yt6xOtsq0XvXFIlbhsMXdp7udZlgS+txLqjPdl/1dTsOgj5mYyROJTSJ
PKRcbLB+jQtyqMflvj5Z52ZBhIwUw03xUy9qnloMSajDWk/S7taL5VaOjnJjL9PR/oLIeLmm/U7d
EKYJjEIThZKSFVeUED6jIA6M4nO1/blbEiJ0cNCGDR8m0wzhQxe/Y5jpim2Prro9kqiqRGa2cMLL
hfOxAnB4jw+0Sx4d7f1yQpNA8QMjwGBd8V/seYVjFPboGXxR6+IqccCSp3wEgrVDPnN3JFLEC7sj
QAZR8ECz6jz3s3PCYTAxRpcILkZa0+a9/Ivxu58ecnUuc3SOeiOKuoD66VOZTP9U3x4aJVeRrSFw
9w1Cdt+e1D7PMH+0NnJXVtam5AKESQ25MbPYGr7+P6yArkVxhf9Bz39y4XSEo/BRa+b8SYMKSe1c
NshImWodxW536cPfypoBgs95q/hEopK0EKTFV61zfzr9RdaRTEgLNcFG+1uy8cn76smlXYs+3Pmx
efs2tdLiBiZS4W6I37wi0PVmLVzB5WEeJ0MWedg75Ay4jLNGFO709YydcsfwE4W1dQCvn/Jm7xj3
BjE1/jxDrtP1nXxfdIpxDytRr27npPenF2INaphCy6Ep9UgYNXXSo1P9UTLBjZMIqCfL3LtnXLOq
7IXO1Og6IJjRm1rOXfSFE8KBMF3eJOqpm6Vu9tQfQfRIPKbfH8X7SpGtt1JiXQrdGMwNL52n/tRs
Zwp2yY50Y+qJe3g8IUBTWNz/zGBzYHGtlJDLUVCS5xT367y03eeotLkWZ09h4rSMpMi9wDNdAd6Y
ht68ZMFn2/3vVv9T775TNfUcUVm9QBIMVbcGahZMFewmr/H/pAZY3ZbxINFXnCyjSnbI6mup0vMW
it0poXM3GC/9A5GGxYNPeHHQxdvok7BqVLiObIlFLRdQqfBskJEZ//BM2YftZqV1JMXWwQKV++Jj
Mloi2xJxFEoTREHVJUE0zdpvk9FuDeewkaNiWft/vFd6GyZ4Qq4gn/mh6SMKMIdAsiUS7FF7EtIH
TlFA4aCpVuiooKL5bocnqW1aqC9YSDGxCQfvd6pily8pdg6NCWW291A5jLMNGGmU1VQOHa/s3MPc
Ziak4maHST4WmtVSBlL/qOv7W5KlDYzeq8c1JvLo7zau3YXlW//VevCa6rFiSEaTX7tHX0drahBG
+crFCCoQnzRbBHAFppvmhDAT8fx4yQuA7XR7j7m2KUOiALT/Vt7RUCY4LwXo0nm4O6dtaRz8cmZp
O9DuXPNKP71/wdl4mdF6qEhgHTZfoURp1Z4AfsBvRVk11EPL1wmvsiWfsqR0GY2CZG87CgkTiugW
B0TvSDJYUA3VzGvWawG8MwDCznWI7w2Jcr2PhISwwM8YMVVysUlw9lgMm3M5KToSDt2IOguYKWrl
5jMvlNRWjWehyKM7bKb8yUbQ4cVpcnQ0Ws4p+u72Kf/foYQ0eGc0mW0eoDD16/pOsar2qA5o/cgW
AcYhgOzo/InmyEYvQRpJ/jEP0K1R/1EfFKBE1108vKqkH863Zb4XsQYEqrEqDjIjFWE5JCHzyGW0
ksSpfDONA6MGpPSK/wK+3yamod1LL3Gz6uZl/o19Ez1hEOf7T+xpeWj1XTBfkU7UHDoHuzGtaWYG
YAmXt9GagbIgCsqfKoYJxqHZj+DdrjXtYw29RTWDHyiOpY+WZvksdyUvwgl7UDvR2yTs2RGbZjTO
AnDT05v0SXvqtTYuRH+bU8zryqqNr38Dm9yjDeaxmu3q7lF3cHw5gv8vdhTwuJW6eW2CSeQlBW+a
bHNzr50kwfES6DWlMlBPOuybg3EEI8Fdemi15X/Qga26kiAJsgaChoEvlHae7rthHrISuIwBGlEm
40StlYvqGwA//pUdWcKslKd5D02X20GNo8p4GzbE+tTp5zX1JIgBsACaCenQhQYIIn/xH8e5/alo
wlTZ4CCdhL+2bI1Hu+XNd4wlIBpqcnZUwh6EvDjItC4KGDKFJXk35N9vaheAt9L3UHkGoWxDuinY
U/v7+racMYU5KLjMkLm4uz2gr7pHdyeiC+5a86Q6lCdWIQktn1BfBhT+FLpJcvYlYVwufIIemIhL
gnI13Q2F95w4E0RbtCFWuX7aT2IdI8TkwjfeXn7PnDY6rQL6BOGRPK+yu54H5DmzMzbHPXbnhJhl
BwkkhwDHCIPJMqqT6NIdaE88Fd7Dv7UwgTyiBhzt2fGpoxGl8lRCaQu1KfukQEAbaPAESmLBboHG
o1gNksTEG3HhbgyVTZq0V4hZMaha8eI4LkQZUzH3z6jSnKEEXtqv158ZPa40/vxzBFrwr/bIVkZm
hNHuOr3XYwGhjsdC/KoM8zW4PvdI21NIm85hiurQH+73YD3jPkvQNn4lL/QNyQHLM19b6J4ZCDf3
993BZ33SVfQixECwXAJx+gQvl9g/Iuav1npjVCzTZQtzEYcs4o4VpkfEcWpamfAJb1JvSC8cutPH
z4nL7wGGRXDQGx3n2G4trZa4hIX4uY2beTTOhEmyPlmGcMoUN+HWvZu/MUXhxR5v/msObD0/P9kQ
rxxVtejbHejzNzR76cNim98Y3PWEqEJ3hd7x2Lun+kaKKpPCH7wSSgAlctBy5nAPOfDFQTO7v/L6
AhwoeCR5TgCOwsfKGuiO834gsw3FSafW2B9dmJgpiQeuphHeuj1Yf9FcowGy4ZIS0pfOgGSZgCzB
0Rjl72/yo7D+Y8AgJOcNOPDbacGNEKqkqGthKvsigSbBPVBI30d8QzQgGh/LM+Gf7EAPBJwvUz+e
QchsXmXuuycb7oPbWnBl0kMYssiEqVbfSNKE9pgpnVHBGpf9sL7Uow50ap0W0hvpaL8wqNhvGAZP
KNLMyPDVllerIxuv41kDK+f50+xfUf5vCE4+MRiIfOKD+b7mXCoHKieACtp1ZkPR09yggefy3oce
w3B9menlExmAGdEnjl7wRsE42Ey538h0OJEW+izeQ8nDHNNlsKQmoGCxxSlNuTr421ZdQi+W0xuS
ddHIngjK5MYllljXuv3HvG3YPT7DcEZeFxED31DQSIlhpLcwMoR0Xdlav8YudQ7/V2qEHsYhIET5
YzJ+Tx1mIZIzkg3FVL9mFwv5j9djbW6rPcwx3SFjxdqkAXTm4SFLyBCwkxZ3bEVUxiqfpt3A31BI
81ydSk1btMP2rg+KfsAUG/scWb5VF9Q4uO70gtTh/SMD71g4Uf3krAGzXM17wbNHIyZgjMPWKvg8
jcsJa66K2XgPYmZooqDeMR7OBeJ7SoKGtJCVhGClbsV/rCdjp/fj5e9OeizCvvKeayoh3iQrMsrt
Ng6uH2SIRlU0TPzpd/4Wip2zHD0XRmB3A+5mUqOwIhnkwiKx3/zjxsut7HR0XdWXqh4lB3Rd2FYs
SF59Yfjnyu+byR1TTCx6BJiN7kV5vVAqjSa2ZgzX/CU8vTdBrf0BoRReacCPof2GacgnhmsrWFMW
ExE2laT3O+VwGvbYmgbgSn5faAPWWp1BPkkGRaJX57g0AWsdWyeIAOxQi9M99RzzIzxVq3mx2gY8
I5qdFwsAgf6+6+fglyxNNKskYKW46ujl8zozqfmqO70dnZJzmrfLfs7Rf6qBQXx9INdvCgOlZZxV
uODoY7+5SVZZ+/AgHiKKgG0jq5MmNJwrHSuQkNGKOAOCUcn0mNbMsTXhxP2Oq5qk/32Yr5rKO+V3
61NbKxVhJSA2BDXsZvpo++vD7sn30J669wvA74cADrKoTkTdVBpEx8bvlIXzuOz3tzs4zEW5SvD+
z106cv63aGQenxnQTyyLcOzuJgyeaaaUmrspLFm3kOXSk5I2f9eSin7pJOgF6mWbYkIx031j1Sut
9TsEsWHdECIKN2r2s3LKM+zoxFwUSYSMJchQ8SnCA41Y9Edhtn2mZL3LD9DzrcyNuqeOIH8e3c+d
0JzJiQTXu+7yzsenTNI7qM2FZvitj7Xv8rcvl1KoB63k/U8fib0BRK3Z3DMlHKCC4RQiCPNb6cp/
DlkeHIAYyMRpB1kvFntFh8/8An7Nt5W5UVxFHdxMDRQTeoe/StpwiFcYSgYkzO4wvDjmBP6RWaYr
BoA3dRO6fhZwwfbu0izEUt5y/yGmf6zgo9+CJBhlTd73vypy0f1BydaTaUvj0Clf34sC006FmH13
0utrROUUpbY7TUA+GNhD0Z+3yjRn7pMG6m1ro0yp8my3Ho3iZAv0M33408NRC/vTsdiU8CH9ERho
s4Rk0bg1aTS85fD+Lq1A167+QuQeTvyNG6IEAi0eVRdp13xwk1DjBMWs39u8NMlEAfWJdMojC8Dx
6FLe69aVTVin/Sgwi5Ox/bQacIjFzKuCvaemT/JYiNDPQ5R5zst9yQQ/LFUNPXLAiqcHpOzWUrXr
mV4pGeZ2n+Qn7NL4uFpTvyVxBqsUsN5Hyp4o1rJQ/NOhH+qku/nk2bExOZJM83+oFgBiXO3ivcw1
bKTmuhMPaqqNaf0RnIFRLff1AMwFe+rg9Q2PtY1IkdP1Bw085SpJfgRm8cIgj0aYZfRoy7AZsQse
A6ih0LiIClkatcwZFak7OsisAHCcC8LD/EnHICN2HS3KuPA1YxDDnw2TnsWS7q8NpDre1Cy95KTI
w4s/IH5AxezdGOaTMoX1BAdKd9ja9PfQM7nQ6qqH3wNxJgjBvw/XJra44rI=
`protect end_protected
