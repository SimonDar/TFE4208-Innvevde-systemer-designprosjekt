-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Wa2koIh3q2mZJjFMMCBBHc2mVMyZDOsxJ1dheym9tUeL11n1zirYe6FIoAx1jIDzwz7iV35wtX1p
PDPaZBmwmtKf0BC6IAAZCpoWFIDuCEzMqO6PTzD/InS/H410m71DVJ4cJPTAZlCNDLRuV4QsyXAS
0D80wANlktcFOLsr//wZm89pTxPYlfMkKlL99ihiJdTKPmq1mzvGDnqtlC2tlX/PNDtK8CWSmZPz
8G60e8MvDo8iXt1Fw/SSUBB6xkh3HJaBls8S2LAyresuc0oQ0d6LJ/x878UGqOhemR5f9hCVuTaL
9if6LCCtJUafGbFCzrvzGdmQzsdHwQDuV1KLBw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
zqIGi2lJuwowkWLYty+jMxcRMlSBSLFTKIUjCCXWs4Kl1QF66mstSC2LFYZz0jspD+Vkd36Xk2FZ
NmrKA+t6XRi/2h9/L7EpCP+dNdRqxJB9u3Knmk6JMdxK1K1Hb2Asd0n7TR+6eUfoMgyxWbpYUmT4
Qp4xR3c8p9ggphSv8rH7P4R2Jx72ibnTyx5abvLaHV3UI+Z6LQ2Tr+JIxMSUXZD065tIIOD+W3gs
0/K5BLJ0K+E3lvIYySHjorg5SIhAtLUhUF59ZR8KnbpOXwDbTXMPr5fN+goqN0U+hJi74vKGSPWi
vn4Pm7Irfrgpm51ylVWmqW/jdyPGd0tySXSgmL6oMRBNSBbCaK9Llh/s/CcQNT/puTkiq+2pfwaC
q4g4f2spiCuUXrF+uG3nb0VInG3VejdE5ehvExENsNMEQidvHsoy8pa+Ao+ul3gjzh6ucEA+UwDf
uTlAite2r8BffS2sgU6xUT/nOyMFKsO0Wx62EAT62RdiExQgbP7EU2gmO7lOchilNO/Y0u6gWkXo
3gU658tf/N+XocwcZZ3SNBxIceBsjza9Y4+ew9QmQzCspIqQJ7hTMFZ28bNIYQcI2o7RgdOuoVXo
kQWKqr+uigRn9k0SDM0JtFfgS12O/mJIlJpNzzTuecX8qw3jFI/G57AiyvaI9UIaAiRo19O3fR66
YwQ7b39aVrhmjJnC7tlAX3xjaKwP968JCpFhdNyDZWWrXKpNCy+w6DOQtg6TDrC/+E+B07reuuhc
AH9ua3idUREL/pD+FqAyQW8CoGwWhwFcSMDlkb3bKWCplP5FbbWoBlPK24FqU3Y5uS005WUowQ6n
67UdwwQ4In+Aogst8Y0Rf+UAxdnDDNNLOx8pd0FCoOLxd9NKTUVaSJv77csqoDwLz6K1PkQKDvC1
GlG+x91aqoZ3rckYtC2O2V0qRmuP+V3MAaX75tcTR2etJnPPeiLw7NsHkqEn8zF+MbisN3L7SS/i
/+oPjlSSSrAM+8pcKy0bhKqGvOxy7oflBYXqvZeM/ueFVz9u0opO2Rdgntikwaq59B4hmK1raqQU
DiWjtZ+LEPEi8bR3o8KF9yQj96Z90fI0OkFkYdd8QKPhAe200gbGizaSJXYgYdb7RJXEQkRL66WE
d3NqN+U5mD+6VxYcmqTZewO9/11E+DUaeAW8CJ3Be5OgaiPnTGBeBBGsdPLCPCOvOkI56MsvL/BH
VKXDW1aj5VvcLTuar5EzD1WgFAdcqQ6eMXA4Kg5HUFd5CZjUuEFoEr0EXf2qtUd2CtC4k6qGkJo0
RI0otR/F/x4DWMk+lrI/MTdBI6h3JgJJqjtvhjQZtVVV4eklpesqo3rxndFkhQoeAJy5AiPJ81Kh
xQ1iFQMKMdX4i0rX5FwFOXN65zKyb23uS2bhT66vMf2+/2Bu3VT1fpbLaC34Hf6jfPldLAMpUYq3
x1x+jW4gdZ+5vCIjaXOVLK71BALY5A2kwqp9FfNWOec9BzVxd6XEDVkIRoM4xF64h9p9BiM6aNpI
EtQYyznUDV02POaGqAYwiQoSCPupvCDC1e5QSu/DsoZDkZUJDL9n33pq+h8DpUvtPsFO5AB3QZN5
JdrRD/kPLv7CczXhiWMap68R+99tQTYZfhYesrsIu8DSyrL1yaavPXHPyH/KCk8i6zvaPpMC0O1V
P1R0zFb/Wlfz+bOPiNFG9l+43ZNvjeOpxcosEodK8tvdW5l2Oqz3hMr9PEW1nKiREslt5XJeLIp0
C6BfDM6msj87NKIsnJw+mpdwNnJppKWMlmXYZJYj40mweCNWBJ8iV0ng44ESSQ/iflVBoVbW3Xu+
sXzx8ajDafe97/U4T0Ttwto4NoL2Op6OlSs+oGmp/cqxTVUAg97Q+lsbaNWDpuF0Us6i7OvRaLWa
+qzaahbE55XjSO08suVEIQoEIfbl5JXZXcPQcqinFCYgVXW2mUP4zPxI+3hm9+/Z/t0H3rgaTpaR
Fzbkn9iUpD/9NGpAkYD0SlSEiVJBSJVTHwRLI9Q7X+M0/wkUnRrxHys3vpfr6B+etKCRSiPfFc7e
avMQ+y0yu9s3wlLuxtwbcBuN76kRnbS2oyFNyljPDszHXyNiOLrVlKjvT5DaFwoviXVKrve77G3s
1Sbm4fMDr9hOBE4xX3tcNgix/diRmMdyV2yWk7XFz0R9gCwKh7dXXwEA3/TFcZ5wn7M+N124SHV3
LefaBWHlUcggyfG6URr/bzrH3sWjzO4umtmL2iH5u/11I6UMDmwoQTEodVrf6t62j+DMWobbayrc
o/Xm6Qwcg1tHp0xFeQHJC4MoIKCDR4J2TcwgQBnTfAcoB/nqv7MwtPO/a1N37YjjtBxRDA50DM0M
F/+DNAwFw2PB8fzDYmzqZnIs6XqLdiIYrKCk+Vg3IjOLrHMHa1dQ3NX5DA25z9lKWpkK2RslF0yT
b6HQicbGw3S3mI4AYmkLTX/DajBejTwu/klE4rEli1C1UYuOyAA9PJnN0BrWxKZlIVepP3S9JXoJ
jQBA98gl8Vd0aKnyLpdjHCyHlFmR8/+9XsL57wPevnDlny/+a43eiXm1c0tdGTkxmuV+w/8nJmkK
mMUXW0jiY5TA+dw4Nd/ghaVI440VaQuO65y6r1YmiplHEgp4535WGN2VVXuTWJovSGeeRpQvo3N1
Xee306Q1Ce6Ft/tOXH3TX76qF4KD3FFLt14VJfHOjgd9agzloexkun6U4Kd9pOEVEW49TWdCPDtC
qHq0ncu9Ev3PXeH7nwTcEpqlBY5auqdRObIxvTGRTX3HFyo39vUoKIzkucFi4xAUbqDXWzkjvoy1
DguI3VSmdXDWdxD8fRuOB2Wmw3GXqeEzpShK/UriHOLuUCCZ2rILQ8hawI/VLC8BB3JdctM1E3+C
6QezszNPgt+eqcLmen399xCowtxIGE+CDFS3ev7tVCLaNelf/00eR728RY3MlUjpYPs43sxyjLJl
Z1mcXTEUz0CEZAevqW2RmgToNpu4Sk2iBoV9SYmVMvyvHwKhdUGFZXl4Hg7Zgr7CpkosDY9MYf1/
W/Ga6pW/gwo7xXBfQGqLAY1YCsJtY5NT1It2kv9j7IbiWhyzKUVRJD8meeLsaBsIoN9A1ehPnDa6
H8+VIGySu1HxjEu6xAXt7vKWudrwVqx3KD5/NZapiayIcT+WMRPq1FujPZJtHSra5Qs8bT4lguA9
HiI1Bnb02tOIkS+qmQlXjipahfbWh9ypGiyOY/1zvPfxQopJufUic4SF8m8q1yi5Hf1m7M2+xvXd
zjYWd+SkOdZ3AsE1X0De0uXIIEh6gh7chu/PH3ZlzJho60S8YW3AzwzP3zEtZEdSS070bSn11vjf
90YdaswabPQMyyjc7y8Ip2ucWwfAieRV82tDSe8gTtbAEBIhK+20DQVokKjJY86pqJ2CLZayUBIP
7phTcF/ycEgQ5Ym5awdupwolwVdYfgYB7uAiBToFWwMRfACbgjRUuyy0jGUJIS45wJHw4hNezjsj
C5wQOmNvJzKV6GwRSHN7rkVvd0o10N9BAvWs/yHALRQDKZWjOT7vTe86TwCzcwBgyw2wrc89ZqDQ
/vfNt80B6RUc5ZYmd3TwF2CWWt3lnDNV+5LtbLedlAPoNJOYQxswfxi5gDtmvj893hwsTZPdcchh
rpeFg3iRbEID4aFTSrTwcPb90B7WBK7qLW0noGCekg+HzUOIzeROBpSnLGF+sELwcTDVTCv1AqQY
vhOEsc4y04iP7pxUAiEYx2Wsde3KS3MW2+UjfN++RpjsRdG75XYRdo9Zs6T/LkJ4l0X1UtQWGP7D
BjqiG5SSKESvkr2RI2KEnG2LrbM26Rjnn+U+2w3aZ02DkpWSyJ/SsycMo3F0OsLDp4jna/2wNWAG
XoDNrJ2A2hDMjYCLcrerURWZ1SLHif2oTfbop+54xeuNRT+25fJSZh4uz5W2MG9u20erOuwe6L0N
K/ItbFo03ZFH/yRgyGxGrqg95Fa2+jwVxR0RXxs+oD6s7pzxWYVL/UUydI0gqk+JuW8tLXZAdfV9
TxsMgeDojsjL3AlVP/D9dJL3xcQCqutsIDO64zzB1DdGk7f+A4IadKtMTt+Y8em5FMQaqD9dkBMl
fFPIl8zXvmCufsoz/dt8Gayn7HgxxQVp9Qu+WUPJFpkWMvDKp4joV1SaFSgn/DlBM6OkBicV/Doo
Xxhu7E/KsXoTrXRfSuo9ioYNBz2tOyqjJKdJVGsudDp0gmqZG1JA2yajWSF3eTdn4Tzw6SQHZyWP
XXoAyyKYbk9moSt1CZXh8Wt8lYaUg+NB3fAHyjsDFnxN4ZsYczujlMUqF9ax6fLQSpvPBt13H9zW
91fMeab4Z1KEjvwIGcmSEk74AhTj6EWHBB3yV8CC9j9AbFl88vPt25/TmSc+6FKwiKcuoN08iCtI
c6VLfKWH180f5Vrefanlq6vPtI/xHtRT7NGxaSx5tzvqx8LmHwc4V6OBDCTiKOfHi4CV1KQlr4X5
T81r4y7frZpcjJSng1XFWkggNHrhPClzdaaY5D8VsvXrCElW6pipHBzsszcSCVwo+WB1Nf9atTbv
5xZ3evTl9pzXUIg8EjTDamVNVIcF3HZLTHwssDogCYMBo+rBWlbdT7IuWncz718sUM0TKwEzUC3r
z7hqZi0gbEPkJQ6ds2hCNY+xcMSZN58UHTbCfvwqApoTJZ/9sLUm/a9eni0Ua1fJZJFco1hfPTAd
s2W8fK05myQbesyc8IgZtk3eEwRc9WIPBg8XRZSbORNZgYfuC6tvwhT52EM2yMtB97i/3x9ms8M/
V07n5g1UxlZf32fN5dEpLMx23SQLP40Wq+Ma74Y+eaLoJB2bh2qiAvHycVBqMl8pQJlC6OCoPkbS
75wgGP/jpL5wb/QCsk9qUHN8RtxbL7onXNLrtAhgjCT26GuK4Ko5CSVEdznBHidL0Kv19Jhx7Y7A
kBzR5QPDXppriXDnWh17uv6mqATuq+cVnmujx/QiTntAYZjZx4142Vo5q6iZd4S0SPXTezE/TzbA
fI3gpQO+zHSiqeTWQ4AIdm11504Tx9bs6DiAVnMOtjYisG9+FCkKpGE2RrfOm/7fvM2KC8dd669r
kNd9K6Ce/6la1UJklrZrnoPy6zBzEk1vIugXHpvfUln/hMMGBVREH25nbYGK4zKSf5gm/IVCYsMf
P/dIQssd52vQ3URKSg03RIjYJ3+7GeOOPRVkwL24vAXdZcUg12EIZoqcFsO4uOQPO+B2eTxoM6wD
RC5pZch0P+Z7LtXThNZ+k6V3v2p9Y5LA1Qxjy1hfBEMECeoOpToaGu9dhTl9oQSK3EsZITwY1vUt
oit8sA9Ip+wOTEz8E7VAydikTl6Q7IzrrWYbPEAKyxJtOvS0nFesMxSJm2zUraqEGdctaUHoU/Ov
R6WMfBVeF64IYnlT9vZ9LYoTNhuNF55f19eayyorSgEHjguREA+YiJyoNrAzp3cRruKPy23CBq26
aKRka9EX66HfbUJTrHUBvQlOYeOWJtAOxBmkiKnYsWfhJ9U+Ht5+3AW4MtpbVH0XJ6B7t+abH+Xu
1lwlQQDzOR3Lz+xbGB76I9RKNqmQqYcSvkTGJxJ/UyG+BI6+j+4c5bjyb4G8QGiamLocNW7+Zy5d
XiNLXM8lpwA8rY4NBI8immggSspuUoJhhzftx44tOMxX8VwUBdsVMH0Up/BLNUM4n+OGfpLjCunj
prGK2VI/2vude4vLlAq9HU+fFeeEvf4eXCNexw9y6iYGJJ3QrZ36pokNe/eIElZN+lCNW67jLcLb
ibOxBa7YNGOnP3Xzw5WscMfuavpF/r9JNddeOdajL4u8ZbvLIg1TsSvQvUIOkGQs4r+2RDvwGcvr
AlUGaaS/mp/BBc/wp4oBEJrWerh2Zo2rrVcEZmDDznvL1oOlZubOPCPHCt9Js93Yw4O1CoRhI5ne
WafdZ3ewe8HNB4MpLLYsQ7BMlw6T5O7ihM3ll1vY3NYOryXhq9y3AMU4GHeMiwIHLIheO2/LnzoP
4tZ+lqlZSlOe+XuMdcPat/TvTAXctv4Y56JZxk802didI5xBIWz7du4CQi1wRGZx+CKgwUEouYGG
2LNOujS/1si9SwbirPZSsmEoPoTzpnZZKGyv1oXGAUvVvbKSeZsQ05N9B2NJ7aOACU11YjYOU0Et
xUz9H0VWKQ4X8bNxcLngu6jMhaQRhdvvwC5QlobQjtSeFn6gUF1dvQeL2iRON03c13m5v+jXKeVy
L2ac/3BDxzIZrGhC+bZpDENsEup4MZwUkAprS3R9TYiDTp6gOxQEXYE6KEJtZqm5GoXup5NxETOQ
LDP2yC6HeQIi5VW95YQflvAyHWUdVtLKmLh/DDxqpeIPKJyjqjiWT3we+e62So+/kdgvfsTrh/SM
5EME7ff/3rPHKYP2uuI6iTzP2MNftcZ8sHUoUWhi+yka2KKmhgVUGrj0k3vI4gq88sSMlw5YJAzb
7bODwEfTnZdarAAFwN1FHAxBMYk4eR9S8BpcJjJ4ZVchpAkgMK+xCh4Pr3TO3iC3GEfNBl1xVWkk
q3wsEFfKQSmtxW03457ZHk1XOU/IXRPJVJThkgG861XJuKjIWVdv2UeJNKCHTYPfw1z0bhOwkzXm
ypKi5UCJgkdkGwLTrGwo5fkQhoc2Lc/91YJKrrut4N0C875yUxcevXlA5tq9hCsvLlz1p7yNeoP/
RiHTw/CrZiYFlhBmH3P3MKr+ShEW8ITmtj3svSXSIIIjC4Bv7tjvLn4uG/8wW7GzysCFfWGsb+Ln
2FsZjby5t9IXNhYtTSq13CHMF1ck7iThm937gkhYsI3P/ILiiX+VER5yFE5uDeqSBZetELkyzFV2
oRQSrYEI5xjqB2ChzM+W0cSQ65vDGd34mygvkj3R0ShgrfUk+zLiXbtZDUB8ePLGtvrWh8onOL0P
LQz/NwAKEgnp9IQaP51icpwlTt14N5dLekV8q+1QN72Sq18XuSi9r3uZmp0JPhx5OjXwB+WARDgw
3wEL5hMo7YHXxrgqsvE6l/iJRxA5LbxVCz+tK8/wIXNyg0m8mRl/dVUoV/KHVUYuYMyIsapIYldD
TUCTeOHQF42VnnrrrBrXqRY4/l1Y0HEsg8+KfI47+0y+z2mLZKsFkjFPqxpUyAn9XWWsNHY1iklt
N4BBlW8f4zJu/gU6AjkWD/u7vLfeajD0+NfXSXCpmo+HMnYy2rxsqXxVCwhSuLsVOAUFFUV3g184
crV+A81e7JLU5E0yVJqJor7LUftVy+wVR2BN38ob4/MHFwanYijvm30xFxs9MW3li2jxcpv/2UZG
cATOrt/K7F94h5jhX7OOoFkUaYQ1u17MyOSqE2vZRdlCdwAK54EzUx8TNvjaPE3fRr/N9YzUBq2A
OnwaLLEAZ2Dg6AJ3tQoOKmR7kotKhOaXpcAH5zvHe0Awyt/zYxDKCeXkuHKLiUo9HGIR+U02rJee
nQhNlgCA7qUpVADLJpCrrmw8TMj7Lm2xclmYS9PsNY9gJVgvgFsjx0MpPcVjn446Z4iZYC542o4Z
Okm2rINrl12cSut+WhD0MyV+Pf66+l/gOzG95lzmeDtu6iq3DDbLSaVirr/ySLz83q7+C7QFP+5j
6tRYGv3aqAHsZ2NOqj3HvBHfvJbX6FB6VfQ8wWO7PJ04QcjP3VtDAXSeEgd012wzIoQUfjnsLyih
NDuLohJ2IAJ83xdQtOUwY9ZBBRiCxIwwwLsXDInkS7rIDk8e8wph2uCF1jy0F/n0PjEQ+tpNalOp
Lo0ASo4LjWgP+V0sP9W1a/zW/oWmTFrumBCffPQsAtO+HbMFuoqtV9iR678yG49cm3gAc81M3HNP
FyIGQuiXKt4RLzBLiH9L38LTvz2Q2J6loPnQZ+A4Oq4M8pnY3YWorVhic2TWzFHz9zq73K+6LEqH
a3xuDIrVgeDmfy5xk1SfRw4jDv1686HGUyENyhjKdl2p8r2MufhV3ZTWJLdBiEXycCxe6lymjd2V
yU8Wi+g1nAiFR4dZ/jDnODOagZLA/rPGfALpxh0uiLHJtHu0JfJud2abtJWUA1qWpknJCH1s1bF9
MVWcwDh8YiULqwVWtkySfAz8c4v84zwMtTzSX+BnkXM+rp6yRIjsgzw8FZZHN+qGSZU+/tYUhC7f
f+EolJyJ1IDMAWdynr66mV76yCWONd/bSHF2hA1GGp7y3tvpu9WFqNVaM1gk9zzzW+EafTl6gPOf
KNZRQuV+BE53baFXN0LKDCW43AFVDLUJyvLIv9JeC/4He5qcditMM/9+5P72/QnP5821C0IZrSOp
CzD+Zj26kYMRcjj0ImnrWsOKTIr5f2DYfUg3U9gyT1Itx4+jY+0pDR2wDNHv9JhkUXmhSQ6A8/fH
Nx+2ESEuX+S1OG42QllQjXFx35NEPH+oPTjWZNyZaWQeS62y2HqtLDo/M+wRcnoOBZEFiV0X067U
XxpFwjsrXQBo8HE23Fyg0Esb/wLZ4b0XkFPSd8c5Hxv/IiEbgf3e0vjCJY3n3Pg1DbfCjF5ort9+
0kNccHCJ1+skXUIJFVwAEOI/ztddfnsLYtdmdO4/S3+gEuM7l5I2rIbmVQwtrOh8IOgKfbpHaAXg
n0ewJKdz8l6rmu4B/nf+R3nkGoD3o7M5rfK2ht+ZV05wx34/WIf8liWOj6+AfSCNpYntUiYIi4qh
B4fzrVsHMLGZrfQH1cP64pqyAyElyaZTAjkNanf39h0UJthLfoOoKg57btOP05IiAJO3ozjIJUEJ
0nHHnqJXehK7s8mlgEklX+4ftZFHwNH8aueoACw3hKRbSJXq81uV2q2HpKtZQML29UqOxBy5JMr9
zYfGZ2u0fVN/99BqFVO5jU0hKOghuuvGdGcEjfGagGqE5RKodZkELLWeAUFtkMejYaskSOdqsyoM
inil1wlK1T+ayKswFnlAD+2u0PuRGzbAb+I0NoJ0te/ydaKtXBIfHgp/V5TRZN8pnj71RGLGhdBw
iTdOW3V7rURLthJy7KLgPxHkhBc6Ry1gPwYNA4AyiixwSbl4zz/qfiWXKzQghFxRsP3Rvu/61aec
YdBVYSqoeGt8yKAKpBUyuEK9FKBTx9iWWFBndV8Tiy47xNpjxdW3kfK7AfxAiN8yDGnp3z5LZCzM
oOMv8niETIQ3rv8ZZ/vgXpx2kvKtNvEnWPJlwav0+vvJwdhXCwDDFNWZPyAOfog+C1uoRzlGv9im
Lnwum+lr7H+6pq38nOVZtSZPcJHT29pIs5/vu4boWfdUKBXYMzR7Ncyj1d9ckurjyUBH3QjuhRP8
XM/41tieAyjNvvUwlA++YKDqJ9ZZhl09+n/3Xzbei7RXce1n0bO9fJaS+klsSvOQyVH4h0TTKplU
eI96AGO+vwYJaiFzp8wQy7qEerAEOuQS2lw7hIYNzGpOMhPO1hTqWWaHBOv68pVrTHdhmU4mOqXt
IlUCc/xYDXd36M8qXkVP2fmqTV6+W40MbZfa0DQGJzZ/xb0z6WUIH0nxzlVMguDFnCatldYO+rIR
VL4xd2ourz5FaSbvQqdTPcmy1DK5ULM/XJgg/kW3CqAEjjFE5YWp0y/b0h86fE7QT5gBeOGlV9SL
JuiV8eo1jAisczWsok7Xsn+9Mc2phbfK1fJfEBYHNhOy0P0zbf0Z/5sLZJG2yfpPy/U+qa0FPO+L
omekA3lqO8sBiOpOANahDQVj82IkFBU9EBMSiJhrvgtrQ4FxFH+26Kg4N+p5WFxKUbsHG48Gnfr7
RqiwMcPKLiHOFQ9pULAnPK8qqGaK6FyqpWcHZG+B15HgwfZWtCa3xSmPEaJzCBzAz7n8rq00Zme5
IPKrsuYPMVnATF/Z5G7lv8t9j29LkGssZvwAABHQw7yzoOeb3SA/Jd2tpo2Iuuqe7zdeC0oHZcde
LgFYTeDB43ApX3V5QszGuOMFiX30ZWBaYFq0E/E6Fil5GaYug/3xBH9ayvzyxb4oTffZt5yyidZD
mQNLQdMcnzUh6JfQuNkeImHXo6g1NDbnE5vGK1SjNu1SYmn+Jiu6f3sEhsFtjQ7NEmgYU8lapU/K
6z5GvfcJf3CINyPqnFR9MPiC0G+qVjgKLlBvcEhugFZg5meSP/6H8WmRapF/w8QrJZSwmy64ghik
U6RbLnIpOUovr1AP+pYBrjevveTsfQQf5jXPvhgXHdIhvPfxQwYPMVEZl0gK9u+JJU/3nWDzprbW
DVmnlBMJugEb6WW/FzdWCqZqBiT+t5E6bX+SX9v/R65mpf0+7ibC0Rl7A16RfuzwwGy1NtHLfjq1
vLUi7bnH+u0/IccEVbMQYtbzljj+VkEatV+pzZBAmN/lPxmXW5VsLn5moLsJ+uK/xS2i89Xa/IF/
rUYh0TiXTG7iNlKoE3owg/ENYLNjT3R7gmg3V7M9H0KY1hlt8yqFKvqkcMwhGNY/BFiJVMNMBLl5
HrNjimcdCA7aIhkzNNfvI1hb0fZS0AEDcsQ4wsSDw8Sf3idniKdYoUfm8XcRwiCAoV1CPA9eSMp7
/FXPpMwz6S81VKKNXHGm8tLFC38sYl16R9P4Ehij01GYl3jEwj+qM8PrVh1GIXRjpK/aGim14Dh5
tE+J+IKAQO1RgiDGmYg38F9l5l5o5LI/SYt2hsEp/Tae7g7MSWGgdkhfvUeWO7dxNAd7mL70jDR0
3qEa5bJL3mtlbKDyflhy1H2n2Z/8wr7n6PTOO4jtvwWtnzRlyg8FxEtwhcA7XhkiQMGzbzk46hnz
TuiBgvDthu9HDJPT5DgbBg52b6W8XAAZdASag6CYeh1PCojPLbYNiQcZcIuN2naxd9MIxooUcqX9
eaoILhLIE0NtoqN2TkZYapl9+89AXX6raQwuqoDZBAoTmMYRTVJESVuUwFmrd4JGxgohMwkWhQ5a
9BwAXwrGjIJiX/u+qXaGUKsOE+tNqCPRZjmBVGXO0yXf/ZeDHbxy6PM/kKCZTdcJS0a1f5T5owNV
4zJ6Swqrf9aJCmE/CpCIJGWe388Nr0cdtDkfBrxw8Kn3mJyyXEw7a7ofv3KvDTfiuRH0S3yKtmiV
RsxQeX4jaHiOPSIbOFW7SJCa0iGsRXx1RrJE5N6xgHLaT8Gu3gdNSFMDITPNd9t28t72gyXI3xxA
pugYHBhfwNN9pFeTNeJVzMJdKOp9f7tPlnVoCl5j5rLanPqN8h1+AyHfl2yhY3qcXYJrfykmeYlL
GHWSoh5VSpQyHLuLqF0oJWY6ePR5tkn1vMgU27fsg1NcMORKC0Z/uuHvbTjHEsATqV6o2kHvhDOk
n71uRK2vS5efnqQDqzJmo8ICy/xeLPEJVuXXwvYNfxgVUZsFho2PjDqNSoROmamlH1a2B9I2NXze
RbKcYtWwZkAqiOnCzmdXrf5OdSwCm1FAwr4vlmNUk96A8RuslMwnuEd0X9trZAc9epWLkuldIjJY
4XoZzNpVz064MgYsjKVxNmbuOADgjO6KKdWP3laN3TZDbsFwJ30pcrC6VbjcFhyoBlSgngihnm3O
k7tYCHwaQwVlUaC1K9/1ESeRbhbXKQIxgnGlfCs0XwF6ouyy65A/PJxfkAOZtb+aMJ8JKTwvZVXJ
iFaL3xQ2/maYkAkIvQF0dtFIsLYsj6btjDKgRSU+W71o4vo5gFzGXIIs9HYaLl4Mvagqhrq1dr7C
sr2OvOFzlU+Bsq3SmpMFIQtAS6ebnJon191EX1i+MHqbbHNHFqNe7G15wfzUyfgodjGh0+n0NL9S
gLyFKyWkQi7zJOd3ouayr0ORSBNhz2hDYKfpF01xD2E/JwucETSb1yAp+CH7xJEHKu1uoXcKd4HB
m7vbNvBuhLwDOZ6nas3wdlJE5imFBqAmrYcSKAkpkBGygws9MKurMHwEld01f+QDfD6HAP+WdYi6
x/D6jUvcBh1L6hQ4pWexHconkBU5iTU/hADw+bJaHAhgOterRzJXl5n1qGTjf2pdSBU4+LeBZK4p
TYBI3dD6bVd/zY9tyb75F+vlOHLVyu42D/BG8GWhVYJqILPSpCvCqLhTpR46a1IJTT0YxbKSYX78
hLPRxVJs77hud9DvCzNYNpwDWhgPCAnlETpK0BxEujgkZFExm9+8TpZCo/Y1R90PiekqTtJP78mv
2GNLGu3jLltHVeh+wP7JLKX8VuqgOQegaoBfHiLsqJVhKUBEctmHDv67j34E6h/JShgZ7+8Q3ob/
UW+YmpYKUU450+jbvO+gUPRKkh3pSLbzRqnLBJKA9YCc+B2zqKrNJP+ScmDE6WF7wmNQpm9hbELJ
1ikLbeFkLmlFwZwdJcjdYIHWndXapoUwemmxH1eltrOKxrefJQ1YKV2sQzNwWyqA+zbxs864rpW+
oO4yXzo/agmFhQzbSx8Xr40rHgAzYiR1CiOxd2aEp+49sYp47xSwoACCaiWSxKS7XyKJBr2DxxCn
qJIP3ukwWE8U6zD9IE88DHCl8cUeGXYlVeNc9Kvm3wxJgRx8W5LDnPlEHCmlGPIQD8vSmXoeTjik
BXGEIByBwEjkCg0JtI8c1Y1/k3zVWPLFDcAGCZUxbyyl4KI8Wrov2TvYH9QJ2xi8d2vdaQtNbRYA
4OuGOvEGOFRYF3iUWbfsrZ2Q361NfB9E54sRf6j5L/XlI/i2mYUZLpo9VvM/FKJGr7HxVRTZpFif
x/m7/OlP5O/3SiAG3GU/smPUA6i/AT6FIIHO76xaxXNak9SD2mANHa0Yr/xoo6LxKlOh3idoACAa
yA+zXgRog9LqegpODFZdplgDNSouS8VxSppefpNmE/2GJxgfRyQFugJgZmBlxg5LcAftVXDtVUVH
pzlK8uPtV3spVdQzhpQrwtBzCV1Ailqp6MWaugpUvasHn/BqRdVuS/excxRPpLFyE7ILnHlJApnB
ihILGVLwpXRSzMpcrhtU52j6zOgt2OCZokrE4Ekz5fROOXrbgjRWNsQaVUwvoa/KK4yA8gxkYiCf
dhzP5vg7B31cMdNCV6lOK7CnAcRc2XZf4cqkgsfhvYAoGXFMHgprY4VeToZal6U8DZNtewS+ZKjV
ySXj4yKFznib83JrqPbglrG/VvLBFKFr8adR39waAuKCRM4hVZBc9IC2gWcGfD36imhaudoaMibD
l9/ln8IxhhUedsv0LgzXPD2DNopgalcJjDNOZ5xVLmvGrZZP0U68HKW3Lm6YToiSjvrB+EPsgYK3
pRGogIntrXxkMabj3IIeYy211CqAAGqsu3zXKqZG02uMgFuNZEV+/u7D/+mc/hYEMCWUghYvSjLS
C+h0m50M/3nJVrgEoMdoCeH5ibqwpvJbEFGwVvsp6IqKjh4LNhjO+9qnmaiUIcZ45X8I+6oM7X5L
HD6Wz87retZojk4SPbTUalQy7XNhSGFnr4R4tkdWG+M17buUc22etwN6bMDClVe7Q1M57jyHTRFr
WQdJmp7Fwy6BGJuhbdxvPsAjC4ghksRAyo5OMhZpN+h0qyXJaa2lFRcCtSXJSzzfv7w006kT+W40
nAJHKEO+lwJSOEgMhO73ybySBpKPO2okN1z+2TpntPWhGyS9+jQ9BHbRR8ufVzA/XrV1HEtSoODS
BNuSHRLjy4brpzPQkkSWmUG5T3ejJ46R5fb7I+wfSjHfS47lZo9flaGuVNf9aYjIL9ndqF7NlU0A
ic1bGOsvhYadeS3mS/ilQgsE5O2O4nM2mssIjEe8kb2e0Ue8OMgbqHNHtfo3UHpP5Hh5+PGy44NG
uCxhgcg++BTsHMwbvpRYHO5qkZuZvQlbjatF4IoIYkkRflMkypxFVeriFSggPbK0NV3YVeNDq+++
MXTBUYh0qYKV1+VBG6XTcXZmJ5WlArF6LsBraM0CKR4NbIS5WlxYpkl2P6xlM6vUGfAELepea4Vh
pRIFGj1k9TbfpfJ/AwbwQuuI7IVLcBZsT5CKnKrakrqIUiVPSOy8zzNq7VcX7aHlvT3yjGVEc0D1
DzzJHIaDT+w3nQZVxMzUxsyRjs33f6qMJhQuQ7puS7GIbuB21kq25x3NLSxN1ZYPVaZOzaO2sjVw
cVyHxEL2Rzi/rtt+FaVkM4r7EECq9jgCq6i9829WzQdWfj5SkMPV3QVVGOKYJ1Ugg/jOWmhz2SCN
DELb1cLCuu5veX3tR8sM10WZ91JKSLQ7zGgt2UGWgTOpM57S5RnTOvpwbYNTrXFkWeur20J9qQLW
PklAG5CLskZQWD1J1YmFcwKfN0I2k/qQeZ1OrjQ/PTuL9plLN0iThds01KrU+qDJVQvpTE9kCDxp
skoUai+qF5/IlSExd/T0k/+Y83ASVllalsym39g+ZgyiPJgaEL4RTqyf0quU5V/LXV+POT6uzMYD
iHcUSVkbDPhMMMIWLP+do9R+5F4kfUACLeWNkR6mfcRv617hZOUSUNAu+oB4y69DcT9jTCZoX2TQ
tlW1xzRQvTlQSkl1YKXf43SvSuEmeQM1GEId2D/oIR4gWLV8IgxG5iZhDItKoeW0rsvvK9AH2Etu
GczkQSPcGKV36VDF5O8QGgCVvRgTPd4UwhMtGU3hjv8YnrQJ1XchFYCJvngXsHQ6TgdDneGcsrPW
g5X0XCzsQYMls2EKxJLk6FSIiwQ0r0YepvOXu5bR8P7Xq/EnyR7vSXG0vJV5OVxEm5QjP8jgPKdT
Nv4gqn0eOl/NMYAQg2Xu6IgOn4zLcCzxiJCyc+FESKQ0HGlBFgQTa5HxMuooqvdnwZ+w8rIwoIRQ
t9qj5yFRV17Xi6m2S5iJfcczkWfjgVCgA/YVvtN0JZ0LNK5/4bHEpPREmVSbSWX3cgHfUA8/lNpN
EgAtdEd0+8H06jr37D3hCLYod/yFJniuHUGK48f7aLMq/+EsWkejvi88Lejm52SPdm6vRv0uYo+Y
upU1YEIaWlmPJksTbFUPAXu3seInNUWuNmqhh8XXnjtt02nt/Holj9jlCxYc8AGqG4L8OIa0PgGp
XQtw0TcfOsio0zmftaWTYzhEkPZPA36yVAbeqC83MxcV4qmtwHtHzU41QbFK99/Ba+ia35nGf8UF
c/eDl40mM/UU26xuELRqr9AHT/lIpXwBRAlVBn1fVI5CZHxxjBIXvAsh30uti3Q6wARm8Agtz/EK
DaNEyXk+w4d+apO/1R8+5lrJ9Dkrq2q/968eb3j0Dwhd5gTYeICX40bbYsFALPNsC4zRubvWSRTe
LkfhD7bzb8AlrIkbFsjGzQHJX1zOZ84IJj6gXlWbUuY94pemQZwbKXaW+ybdENaEg0PbzO7bF/og
aC44fwYOTALfSt+8isR56A7nTk6tLDo7NtkMn5riO6C435XgajVm470HcJAY7xxpdOnQ29CA1JTG
mxZK+MPdn4TpPzPWsiUg1kIzgn5HbZ3IXbqsxUJbu8bRIhAbbr4wbxpiy38vgIhDOpgjRL2/aXN8
bqKzfwiUy4KoL+tOQl2BHvetuyT3WVwDYH5APi4ic2dOsQgoc7h2My6LklkK8WFQaAFBXTR4V9x3
yqLh1o+BZMvBfwmQOkmGfqd89nUOQFgyjWcRzlaCjc8anJuqM8NCLvwKlCBUHx8LN5eJWWiOM4hn
SvH9LroaOU/E2WooixetlbzhVpf1lFOsKXL5czbQ9/IcHArwDo0dBMeKQWXHaMEvA5RFd45hOgF/
ttsEJilOu/e/8Bd06Ea/hvZSuRcfHb8Tls7w085sLqQGuaqCHIHQOUQZw6aSn6TrOKFgzR+uvca/
FuBalx9XxyjcuLosmS9B7Pet1c7L8ytXT/82xUs3srC41WfoidZ2qkV1sz4s+kdI4WvWa7RLwbRx
30+xxUv1aBYxFLvxKbz+xPsWdQGWO7lUFryFZLSChx/SlgfGAsts+y+P7QiAKegVGlUr97wNXpyX
Nx44nOnAZoV3DrybbgNtkfiqwTjQKakwa1PppEV1FBramgaYy0pdHKsrRomYOeTVole+ceQl3ZvR
hd98luedaYezi1x7E5PkB3yLHHKQJ82+KDCs0AcmgQpd4QKQqGd5dMAkPJbzv1vExMQS385GB9LV
txPfUd98z9m0QAGfscntRWjBaJt4H8THxML235QkSPY8nrIzQ8aCUrDFkq5tUeuQvheR6zxYxCSY
JbhB0K3QbABO4c/diK1e4/TqjM6ZJn/bHk/6ZsbafMtq1IqTool52x4ibg4R/xwV5r/XFGqu0pox
ZS8/AqFQ9uSNClsDhzeIUVn/NaRUrpWe8unkBBaKTM46mIEnqHnQHHzep3yEz/5ptl4wGtxXxYMq
Ym25KFsqxI0MwGk/++BXXW80eHGRFc8S+2/psJaRAlnABmcegMu76RmL5QlNUPoEt4pl7LdhsGZb
Cr0JIXdniDJIzfMufmO0DwkxrtxDGXgKrJyyrWJgtrJxqAwY0/vkIAqfukwxlgqd7ZlSrm1Tz/yU
AkHEHzwEpOtNY4gPQWodNuPReM6DXbk9tsiuJCPtRHUBF6ralCl/P3QX9Km/regvvIZxtjVr8iSY
sm7FnTkEFFTEA+cSvjpQr2DWwEDMufHEIqA9tenacJEwLJEoOVcdXOgwWCQ/dxPwiZWJBnrekYbi
7kwedk4i/zVFNGy4XtHOEfegobbfs7zTuPgCSCQg8XFtWqyh85hT3XxYzt0HUAMENMaRKsVXkUOX
dRGzcOUG5aGwRVhTnLABLknhQBTmzxyYM/zudS88SGk5AJM21vVNsWuGWR0as5LUucuJX5D8NxZM
n/UWtstbRIU0qwZGGjh/cI4ulBNYScwZA0aapc5AVGnxII0G4iR/jKducjUW2Lo6zaB4DX4GJhRD
b/yguLYIVGMivEr8HEUrbBwrxxr69aOf38A9YTw8JwyY3TZ0Ethci7XV8VbDJSArJsGdwbRm+Off
yO9z309Ef7OtJHqGFL4VcK92zcDOAPvMgoUq9Eaz6zDxxFVcre8fQnCQkt0Xp/JbK9tT7AtoUI3U
nuTK+qn6BKERkWyp+NRUfW+GUHidWHXGso2G4Sbfo2iHMllnIPMbpOgDC+0Ezvb5GAm0TMRRo002
JHH+VZn6+r6uUw2UHNyaRlDfXi4SEKmywPpXxXChBPj6c8vXiIVgTLYwUfCo2rE/PYg0+qqW+KvS
r4lLpn4Y3jhki1aQIo9lLATHA3ZIy5o2ORWzrH1F0Rp0VKaW72R7OtbUCKZ5f5Yxw6GNj9wY4tPK
8WdfuhTPK8pNGxRi68AH4YQLrGjuz9Th1W+nfc2vKECF6L/kCQ3/2neXHfrxLG8VX47FhfRrJXRL
aF9uQHERuCHvuPXw9J4INZ0cRBa7BphoTOyiLpdLi3fi+jXD5g6f4KiqShgB5qOvdzaWJjutM3jR
HlfT5428il6reQh7/AELaHK+3sLofnVs8pk8t5cTlinFfNKcOFOUryqRo9uzo4ZqL1Izb+2tw4RA
vApQ+a7ykQLEEi9Gy+0ZXL+eW6BDJOp3iDQCQ4k1AJDvyiI+9JXfw11M92o27iGQzqQ/WS7ixuLG
XqDsurxQHlsm7p0qU8P0CdYtWVFwYqOjdt5iTAOQ48CjXVrhEYZN6nowcxZeM8qfcDCwp0Eby9QB
6NWmE31MIbLnmAwOOsd1G4tTaPXFvePLa04LJ4e3hKgQzVRaAx87IC0sGKzeeNGQCwR0gc9UbelB
nfodUoAeMnU01HzgHmdZ+qqQBrATPXyCGQpX2ffnIvsxiFO5gGKn62LbGY8mBrjpMJDxbJPOE1Rv
GEYfR0p6Pil4wi9z2X2bmysfe/VVBBeVJk3cQDk1eGLxFZTpLaaTAzsuBBvXswtkyBiTZpDHG3R6
aMULTEPg2RsRgUySnK/oiW5qNQDERBgr9WvynYVY4WFzeuUyJVsnqQSRz8/VcpupGG8KVCkCPukC
Vbb2Kcwh3EMR644s5JAwWiw+v3+HNij6fDN6n2wEudIGQ7g7QRjfy+rBEDo6FiCtsOE9DEmUyka5
z+4kB11I6QIVPUjXp6ERDTaCdzSBkeiSsxUfitlJqQsgHTKtDTtLQJatptSKKD65l4sQBz7w3uGu
LG3qyRmqDOUaiaDcdCQDaZ/T4juXJ+yVCrFmZh7Cfm2tp/OHExqpxHaF/VMB4FBBm1cwEvk3Xeqh
40BRz7DCNvQH+oWcQE8SFu1md8FH7HqWwy5s3Dy4kgsS349aDKjxPF58G4JZadcqI8SXRIkFJujI
ikNtyLEUXl5FZiakDzRd0IQxWMI2s0IGJK0sO0DZLyrNs4ltg54tgJyuaWeQPaNpVxeuZHTtbmJ5
FFPqABhSj9TOSzIVGmDcg49Qay1Pe5DfWPm/V7VhT5GOCwoFoELXo9Ferjziovc/uroWAsF3rZRk
E5VXXPdYcmHim0Q+oL8AaNpdG1Zx78hZJCLhVf8+DiWxTFJWiodW0+aAyMeI8oyf1zfDKED+NvRb
8Ryzq2psgMfI/Asegr7X7+GvZmc+P4tmI2JafFDHrKL7FSldl3+fSO7okwq1tW97N9iDJkk//VZk
4zfQVZBcK2e4xJ55pMtonGxabg8FexzikLMRrPs++76uq7mTRef1ma04V2JfF7G2yvGzSguKNgRu
IwHEwkV4t/LjtY2uEpGbNfo9bQQIv/j/uG90eX3VVpUEx8wZ0wUfyBnHDrds4p/r9gysrQ4QXhX7
XeO/AcRYpPqLY6F0jx39HkI4UvyU2XdZudVpG0JKma+emtTwxO6zA6o1BBwwZoK0QJRVnth3f6n4
y7Xtl7ODksBsM+FBnL+B2zkZXJ5kE9sEjbd+AHRHm0nR5gtcyj+KCu0ws8Pf4Ro89iqxAG4NPEjg
N0hjuBTMLCa+MLe8vgnbpcJgdAZ+fYuErKmodNH5EukGr0M9mVwhqCbFzxQgcmkkn+qeNQi4dE0J
siwUUZ1gL4mFpHKpla+FWzqR+EnPSgGRB3QW9mQPRaw5np+ax6yX5QJcPBnXjTTx9VUiSNA8em9Q
wwwzaPwYQG99wzffkPM4UVoW8v+lwFFokM5jqq/Fucxr4vAclm20LoWNsU4EFAHTxnP1NCF8YoAG
J757Drsr/Ryo/zal0Xg8xuySwZPymWKpIamegdwhNP6WI04XVMSZVe7YRUXXxLWkFZFmH8zdchbE
yNUpuC03x5ZDAfpVnJj/u1S3YmuGbM3kFHiADGu3EX5tVRnOCHLCNqmSU+jhjI6usPPM5bSqKlY3
vLFPo8aQ98VNuDLe2AFGnYX+ld86C1/J7Z7DYEyfWn9oV6q9bEcRR2X7P2vq2/a+2RiYbnNrJhDY
0UNs2RcvFu1ifb6uPaMbzaQYJjiuOriFwipIfwavfozSE/bHyK935AH8gR1hhArjutPjbr305Zd1
/SqefzwI3plqIvrUKqCD1KuSuZSfBwgE8UlNiKpOtDRiXOlCCTXffDxA81uWbxpqO69aU14BBdmK
rorAd60i/1tdPGz2YdDYiaeyC01ejwrckiKiiidm5WHYQqpm80Ry+kM4FSzCAbcGlp3IPEgs3tiN
rLvgKX5P3r8/RIK5DgaQFg4ethb503YOWCVGfAYpCDxaTUJCAYaDF764hkikdfTMFNXbRzPWrhEz
9xaqdXhx0mjlQy6pUo/L/1kLsq8p64FD+PZo06eLZx307p6QDC7GLkM+Xm3H+YdSLdbNIPLJkbh/
JgaZ5I41u2w0EgGj0manjFkWG2WG+Jwty8OXoYT87fdFr0dTXwLbJE8P+ZCxroQ/k94Y1T/Cz7FD
gwGzt98Tz0GpqWWzCZwC709QT++YnV6My0Agi6MosY4vavM5K8wgDqztonyS+Untt+RRaLS12nqD
+xzoRRq+JmqiQWvI78pIfho28y9NfiXhaT9fQs3WIs5rtsYVfJbNpVk69yPNMRqWTMjlZp4Jq/l+
J7l90bgPjE2Ln+u6XupPj6LvdXsOVkmlPTguCPlE/1QrKsQ53tnozzW7r9C9MMPz2tYvHv3Pszr3
JHwSQq1DkFDBI3A0PKupCw41qLH6nCYGx0UyUwH8TxgrLq+Q+pjIrwAV3zWt3NyrCJmNZ4XZnu5n
ndjMQfR/nXXts9cDGO2sKRV3EjP4P2IpW5JNhY0A4sSoElcLD6jCmWsG3cflY+SvlPge0EpRqFST
DMXh5P3b/tiIKGRdEABPyx8guVbrti199xoxbF14BkVSwDour6hMtDHOjo9i5s7UYLAsmSeW9D7x
k+j/2pPEh1nkE2ZGFxMiUuM9+/YZmtD9w96ozLyZfCV5meeF7wGz1d4fEb2RCKhdP6Yvptyn31Mv
pYIXuDNax1H2jQeEkKLCOp/27eMVLQaJ0B3SkjLD6pga/5qAMia4PImUFlir3KfE/icJB7QBjVi5
QPfzfzTq/P7j0Z8e7XmJv7fMxneHCiVxjPjlZ0/Da5W8Zwuan+xHRnmKRTlrnSt6Gp34I1/m3ROh
dktyeSMH+LwSQj4Kun2jffElmeGRc7GGyOlf5JLr1wXCuFa5KY2NeARQBnnZEareZnA2Qg8M65rL
vdOOlZzmcIgsu66C3pvWdgfoF9FOly+3oPeX3rCPsO5bW17OarqeZdTp8qnPX+i2nlsGUxUuAeh7
l+00+cdu927Y1Zg0uORQsNiju72yCRh0JsAJnfQmwViIksvq/GwmacCVMo7YT5rHZEKkm4KpW67p
RSTWTA7qx7SoOgcgNbUWI0wUqXdCcb7GhU4UqbGYUs+rcTs+3Rt776+d4TjRyh2CBxp1HSA3ewDu
EgoSu03wHWUtVs15mTBiABA9j5yBtv85/Tj6WYHOKwpsOiYsYdZITCyLdFxM327FSXSrsPyXSEby
bYquZSzH6VNp3jwIzDejTWIbUYNp071869ZYBYXXEBLNKXD9Jxve+tu75/2YYeWC+WNty+ZYnmN2
8fTtPbEJkzbqQnX6M8O3Y+Z2qHPOBCRiYPP1xcxNbzVo9XASWT6D1tZKabXuTYt/Ae4DH+OvS9FN
OReEfrRF3Rr6ldxRGbbchuWRReiJSFWCANO/t29CLxak9mQWzayf4+Csu62fKN2AXUUCX4dkRSgt
Nisw6PlY5eFTv+ykKIvyh/ZzHQgGqD0wuMPg4/2fzfIMxq/TYOGaKIjgD1unHOBgv3uLy8XmPkDq
8uxUWj83k/bXdAXAsV78BJWBDqwGGbIM64/8SDvk/s2LbBv7yR9P4pirGk5BJANppngwSb82qOD3
popoJLXFvn4h9cEMX94ASxp3tVEVIwllnTZYUyf1Q/zboBa58cnu1CqMWDztsVlpmqCIkWNdnEAm
RSHV91/iK72Z+CvPBrA/Zb3xqpBYaUFavqlrMAwE0cgAXjObTjSbgyCbbLnXAQoEEBeXb+N1wFix
LwrPQMEYSp2p1/s4cJ3WBrJCmwDsSAW07R2WbzWCBkLeY8wxJIhShMJfnnz73sxM3TfSf/b5eryp
3XKvs5p3npY5a5gKsVcPL2gxRNsALr0k7/Nbo8/Vv563LRa76GvZmv/AcTyiggLFuAjgkp2XJo32
3zRW/03wRw4Lsw/u1Rxn0M5mB99edFrnupBqVh9YSEhM1KavWrg/BzpHt9Df9qB+pb0+dMCWHw28
dQydNWsm/DIh5k9mNcFSsj9OlvXcsmkFouFomaP9GPsCyw2jXlOa9PpGPQKO0n8AifR+P9gon13m
CtB+v0C4VWYKvKh3uUm2zuWy7saqkbRB+ql8ziMWo1uY9PGFkq0zmNJYsNfwXEKiGtfXSOrBu+/+
qZzTMkW0/45f4DZrXlChiVcxjRf2iHUc6vRIsRy+LDg9Fw/1YJg1NpPBmqNpyFn3OkDJzZH4bwXh
3Qbsz1YZ+/hHTuNORFjv6yXaQLANrtdl0am7jA0JdPJfKqZqkFu4jbUzQvVW8Eo9MGBUHPHmF4iA
wJ6kdhXeMpA63yHDaS383jHLr8DqaeSU7kQRN2e3263VgZ9RMY3zl8SQeVWKZjo25QvYT3nSCTeL
d5LQhgdoIzqZPuHgu8sOqwQQwn/6PtSn1i2MYV3Ay9jNQQ5FL9D2OTokI1B3kExZLCW9nDXg1cCr
3aiI6k/JFqJJDaqfiKPJ0IuFC/6f1+GY1BQ15APA23Ix/gwPjEhB9RMkv/13DiOFkHuJXc/hb8zd
jJWk84NQsIs0AOTZ0IKCGzdzyYv4f4m4K/X7zi9a5WHngv8Ch1JRWF6LpuP6wL4UJIUEHo2sCc7A
6ZzlZ5UraA6wiCcmqNk2Qt1hT6ABX8p9U6Prk/x4jsDnkv0C30893crSPj0+IJBi+ocUup2JvN2/
P4kLS1bbCk2nbk8iSrjXG3IbyPKnvIk9wysTlzBDe1lG811Z+GIBN5h/kT8fOv9LbjYPRioiEVA+
tYI+vsFbqqhuvGe4rwPhHCEnjIiKEVsj9C3L3EG1RW2nzwy7Jmpnl8IPrb8LKld0Ol0MdOqujNhN
W4Cqoz2JI1uTYbFubJnsmYH9TJRNbyK/0QLkXLt2cDSCL3mWZKI8UcwBLsufxQzYfkD02voN3I50
IvtGMyXabQ3+5jQICgiYddXdSoG2GVKrYcLrpdd+ugY+E+pcK2VY3u8qKOFv8F7rFboIYhtM50FU
n5o/73F2tbBayR50RPAWthYpWICywqIrT1HKz9rcjQO7pXTnebpcELZDtcwo+hBQJJsPoWgMl3El
KPnZ7Q9DSf2UdqZjp1/q4qfwWRAod3eY6E6E/j8rmIDang7EGnzOUCGQcpHJgIw15pkUhNnmiIEn
JrluY2KFNVIJMQPRReoUoLlPCz6Ys9UkaPO1obEHtgc8BbujtmHEZrRuIUJn/d972XKl/+N6a3Qd
LJ+n7RTu+jlqF+EvBI9pXYG17WAFFiFVszPEZSE007IshZCEXA98flFxP+EGrNbVEX051yTZlSJE
e7tc4hEDhmUjllA2Tpl8brhKtIL/VLOlKEuDvmo/5HqfxVUFUKKPGryBN3JKZz0b3y1FHeGV0fpZ
4t3EBPZxUsFblSJhXnLAmqzXwGGUpJto/I9p0ArAowWiIcLFMUy4b1oMU7m4sj12xXbyyAQsc15B
mb60bcF9J5WODTyU+j0quAAQg4d6az1wyKuNfFRjGjfzZqXQK+z7bXynr3DnngSHWbzyOW56VcuM
0e0eL4Ew+NsjkMuMECzYprJlgoaDnskjf60AzOqICiAcmkmfdo7/uPfCiL7WPiicUOK2Y8o8kHy8
Sfcr317jtpy0I+MA4hSCd+ZVSKLzSiP3h63iSFM+r5+uYB4juz5/AWK2zQmxxzeNzSc97vQcQiAJ
RxL75XZLBy/ByXBTfK2uv+g5FcZgDYojoUbL55lMnYsuneuFEt66EdmjD3OCLgPnvMlBN/EpaqBd
tweb1XBuvnaz/sl05Gl7leGE3cc5Mb1ixuOMsliIQXV/mN3GZ+RIDPzmshrxZEiD84DHfk0fRYIO
4lEQSXXcRFCLVy8bXIAkfyxZYdg//dJZLktv/ldCExECgzKEvaSALPthw790E5tTlsiBfSOeOOpX
nVpTHrCdqXruW3c/QAS0gwPVzcLj8HLcTkddgJwtjPVsvzTYqrsfk7gN1p9IWeJiutk62fV899Oe
NQyjAn4fBzoIAvjQyldFtCHW7IKRbHVTAZTWScJN9v/5fuIdIMX48s20qQqm2SAmHFqyAcb5rwGx
5yRm/c8UhqwMBbUpi5oZiqeLh6Cmjq9xB1t/a82Ghty1MKHzMvrwSMbffNvQaNSjmogM8I9/X+IJ
v73TtmXV7ISXgg4IWjGSyvlZ5bXE8AEFiqJhuSHIWk/OCwFZ8jePWyJTp4VUT3qJgylpmkyW+LT1
CGzM/aPapxBOxyLK9VDbC8c4QKca5epRVlQycWCeHPVmF2l0Am3eLglpEoakORDWFAS2JymbDzAB
Qzrf/mD3A3JqheeYDhb8OFodtUtNuIFgvLersbAGPvCbnYKx/3f396174SmtwiX/jseKNxU++fyk
DL0rGmepESV7BvqNkjDG1nlly50iHBvGVEh6ZwkB8ms4vjKecqcQqfaQZHDTgNz38xtMWjwkJe67
77JKglcjO6Y66Wb7E0k9g9psD/T2nNXSwG6sJxbp13xJj61QrEnXlJ1epsQIsMI66MNt4CFh0BMM
krKj117TZ0wxGeVSZdrMySlKBStuiMekC1pqOkqKuJNI9jqANgnOZSW/eGjrdoiD5S/2mt250hWk
mUgmrXLzL+DJjM4EkhW6n1B+GYIDz/5vd/8jMRE+O9QC7RLzxhdWzaDkOyPfUYWPe+8sQLe2vmru
8En/ZJoAbub18pFG2k1TnLd7G/UmOULtT6yOHAWlnfqDJOBNhGlJgrOPs5XKkpIv1/zKrnzLeUtu
dSo86OfoAmRo6wrdKRkepwnYFVwITsG0XbaeKYwzYrQZJ1MiaYj7i+2nhwyw0Ue/0b+9PI8nc8OT
z39dY1+HLsYRXeHktXtGQ1dW6+d0HyM7oAf5Nw9tWlMVafqXxAEz6io7wadPnmPnavS9ASwYwmRo
ClfbaRc//aDMYieYarD5vUXZKhiEuIgUua5AqgYqRMV2+gnGKklNr/PKKTW8rSEIn63X33HCsYbl
3vxuILg0/awc4CDfrnmpXu3Hbyj9dR+UuPxp729esYgpGHKfMUwep2/JFyadGuasvvnjQGZ1mABc
+c1Lit2q0zExwyTR9yL1hVdCf2SnMZf5cfV9E1NYSFVDZt+jDfFffDGozB2KdBTOB2rQdD+1k/BL
3Sx67N2f9DvMS0wv1oWtkShw/qvEXC3k+st+ExjPE091eXzlItrlergpNeFbmarQgVYKJImmbNR/
8Lit0jBcPJ6Q9PVNtBAF/7ZrqDR/Hi1pdmkpe7KbZIF42ER6HZV9jneGVzJ4z+88TVrlrV1oZC4p
mMb0S/b3R1dmd7T/eZbc66snXMPAquX9XwmNcNnY5mPM5J5pb3J9iT2x6ARjGEcdhqv+0+BD9T6S
a0UyAOu3UVj9jCIUdON6YhNvIJ53EJgoAnoEUZXVLVD5uTPClyFdUwXRukZWXE5tv2lORQInf+4j
bY2lh7I5fTj9i69TW3Vw9QjPVWeCWXJTkNfE1chc0C1w/45tnKHjiep/LXLQ0LQWOFo7J84VClyS
Kw5kRRpdLd/TwMVxyzJ0LJ5QqTWneqOs/ZkU1byJKaZG+9Q4LFvXh8yryoibU7eZmaA/DC50h53z
HLWsV+QykxbjZzIMEgmMgvOej69Ag9TZEcb3Klhz2BTN04rHwHzzKThZqFhn0nMEd6Oyjp6tVIpQ
4FgJPEYFqMvlFDuyuwXwGk/y82mK0WnDtFugz078w4kDkwCgeUj7PZU5T1xmxh7HlV7G+xfJmRig
Vt3hnLqmiXheeFc/pt5/vzk5h23c92yvvHo1ME/LsdSSj71n2mTcb63q9IuVePGqUWJSRC912qym
B2lqRZ040LGOmRhSvruxRf9PtzH27rOfa9FNbIVkm7f974ikQga80zaUjJ8q79dosMQpnWui+s0z
6R6Ih32O+Dbmc6YloDYRdFNFs/+hhzGkiWAVeZWm3cA+eJ94pFgZNVmTxVPOJzkPtzQfSPrxLdoa
Fr6Vx3BY+tyHFhNoDKobRFMUF+EoB4JA48ICvltYXeP+uoykbXu8cNGyxy/IAA7NDIGxK+/gSobR
HQY8eKDToEJBQHXiyRwM5ibmA02K0gCZWC/YWYdFXk7n4jAJOEulMkSi1F6rRctm/Dsds2xTzqQT
ZtSwnDGuI7ZW40X88XIlAeY5QudbwJW5/C7MrAmlTK/vI9EFDLG3iY4o1iUcCmG8xXE3xOXMt+UR
RxnkrhIlMCE6Pe7gVyJHF3unzAZy6MOTAUV5LUPOmx01vKRQ8HBZ/pgb8EbwAtAo6wDlBNVJo8Dp
WDDWD4cmbRcpbnCnJwBi+smPSCrzsV0eNO6+AIT9sfcIZVNelMN5wR7IJNQRwn6Qx5hP/oTataNA
lftTi/iatVi6Os97XOo4C6N/gH0mwf68FVM76WHM3RC3gogEgwyQDWy7kYnx3w7LNS1TM1Lf4cHT
EOWDAv0QtapPvmzK6ZDXQOQErKt+XHqZXVwds3dy7iRANfBYyTDyRhKKFgqeT59svOlv9g/bq4b8
hzQfBtuSBPwQM6Ka02kFshlcFS+XA7P/R23Ch0Nxq48xqiuycrkNHAxPrxSC1AOU2sQDPzeGjQ0m
wyPis/tVbZi2eIyAiylPT4so6QDTSm7NBFEFZ4TLLIZfLCvvuMu3fpJ4lTWUxf3lNoD5jJPOE8WO
WCEGXCuXoOwKcoHAcZGZUwG+47C+BZGSAL7MlzdNsAdle9CY+11g2qWD15UFahf4/BLol5F/ho6D
v1Qw9w9Jf/qFep3IPA60cEIA1Eg66QCYntuOYVMkqZuNJRH64xBPHulJVjRGeNQNvob44vi9EkIb
i8vtXWqi0+iS9yPlSr1kPQ/kZIWNgWpqbgmB6SjsYisBe7QeyCZknbwD27j6JSM23tVspDpD5LIJ
T8rPqdQIW9SKnMejaqBXKVn2fAAxB52OEiU0R/A1BYkvVw4y0A2tNvcGp7iYbRcfM6R3rqUZCafg
rf7Wa6K3gz4KOSCFGpGmVLd1n7pTBllgT6VmbTv+NHs3UMVHuxqbS1vTfcxICqtR08g8WUpd5MZr
AGNZbeCSMJctYpmf7MQTGCAs3q90x/fZkJ0dd6W5dFmpj6kuBgPqYZvhAi9tD/aCKt2sJFl5Y7ET
wLDBLpFry5pFMWw5GhoyfOhNdzFRIJ1a8DKrx1WgF+OH8UV5sOh9R9flzTGLx8bRVWIGeft6uFBw
tqRNsX3CiBWZhlHiPqufeFwaaqlvsbaNjkU6SR0jYQ6dVag+r4mV2OLyX7/3RiOZulwLB1r+cqQd
rl1AZF6XRLzTNtv6znRq+5q3u06vMxLzqYdlA7CF3/1qFnnVsDJWn4EVTD2d6UhuFPhr7Ni35e8u
sGFdDCk+n2kM+Ck8pKZT22XRgrtrSuhW6T9InWnAl1FUyVAVcjTIVirgWEWjBIzmvzofG+iQ63Rd
v2K8M4ldQkckjTOQyzeVIcxvbVLDfUnMwghxxiIttJpUcxZvGaeOJ/19jQyZB9p+ux2IGQqO7aje
42Mye9azPj9q290RHj1K0EzVW27J4JU2wOt3kv0ESMRSr9EHBJ4KduOjuQ8xi24gy25wHtSwjYdn
IspPlRzgE6Dc8P+ar6ESakNZmpOvextBc3llHUBpPk2sDvgOEbO5q0Vz8tY1LBN9fpucsUFlA8iO
jYIZf/djj+z/QBEZhJvQVzqWWQpWqcLKHcB20BBNk9uRRIiflhNwPER7IGl7N1hFfpsjxHlPbHS/
asTNdZ54JxXUWMCphcFrHV3OvNixB1Zg9EMR+9/MfYxYw/ib0nQYFHhoT7D4+Pjj05jEfIZiZwWE
hNT2/EVYqpDEnZS/xWJIZecxOfw8+0O5f5Kf55Yv3rqIbGZhOO61TTcuT2pNvc/v451sFOObphr2
vCpXwR8EtAMx2aABx6iFtI44R3QqutQICDa9plpFO0c1PMv2WUA+Mv9tEDbgfjOIhUBJmAg3YtCR
hU4O2+9BF9lf2mqIYxCMyGYbGcptZRbiLUrF08LlAbIGfBaffzcqFepfxsmrVz/gaFBMfqZWJnjb
sXP4f0cky3Gt9LTStMK+Dkznx0+N3ke2fMZanuAg+EK8fVpvfJHDoO5nNnlcVIyAq8eOh0iHWTMm
7uBo3iWIOwkyQJTzVjAs2bQjCphCYCM9G4QPCAi5bf0dtDb4yrDtiMtFoGWs7xNHEwnYft1yJjz0
SznCTe6X9/NtySwo0mFRM41nM5lG4r5s/8/YxMRe5Qk5/8YEEPlYS4uAC3cT2Oy+f0xt25wxZTO4
VfEiB9ulDpAZfkmnc1DXFQaRxjWPaxEipw/DyMneuMEW4KzMAszdFrzeo0oqSH6b7sVwkwkcMILV
67QSVCrqUTF2cEAPV4vH27dJaJe1yV6FpKqMdVmxsLFoXASDoTtxBBC+CYYCKnH08Lmg0tAI9XjE
xCv/qtzh9EvfC1EoyVez2kyq7+Lux/9bXlWj7S1x+J/Kal2ivhRyb40QvBQ3P0UIqeP0d9OQjVjY
BggsHedim9cDK52JAMf+nU+krljhqzyXL2o2VRMxpGObf0CyBksbVjuRxT62ilHpDGj23otQpUXe
O/d0hHsdcVR4SgF0JCdJmFQXfW3q0kASYd6oSNYcWxZVyB/kDcGPcC9KGhEynq1danggixQyR0lY
RHrkowbWMdWqeV6r5h2WOWSuH8Q0NqoPzw58IfViJvYgp57Q11CROydml9z36nBYzK1oUcOMx96R
A/QNoNXYa3KOxHH6lX5MBWRh587uV4UiXH/O6zYxLbFaNJhcFnJzto7/o+eJWa5FBE5y2gOGy7Oy
SAXB50OpyQ2LHLai4hRpulMTM07FIhnrqvxSCXjcM+YyZitCS00qpxo55BAbCEhJUFWFlYY2iDzX
PTwqhA5Rjmk2675Q2cS11gnGmYF2wgpIGyM3FzOysVszCt3YNpI0ZzvKfjb2zNbbiJzAcJrGzEiC
7ViTYZZBZ040wO1hNYGIvW/iaQ4pml83lJCHOIFIL+5gTc8NC8+Id6Llpq2BnxyTXoH9TYeCjkSe
GtbODzWS/S0FIidhdAwonOSaBqjd6gA7FwS2yEk+K4pKC1BqRbVfPY57abl+vcFtD+bhAA6HJeCU
01WC/jzpa6kTS03j1G9nPYBs2vsv6mm8/8HeT7+KgH3kUqnwIjM7sRb8Q0QioxZYlAdNVJWGeNBG
R0tQGFqmN1BRQhWcZfd7kx1v/Qg4+1lGrWoGb0Bsp1kSiyDFM5R7hxcNlL+/A7czTjOdNhV08795
9U3mRX4MyIt7jbagVZrYai5KJ/+DgF/D4GlG7VNXMc0TWi25O/p3DpRn+1/594+wgfPMJ3s6HBvl
uy8XBJtijpPAYHGAeM0et6k9QgO0+o51oWitLjzZvdScqdFnmadlwDOUl32rhGMkYWIoHRqhRK++
gbAbfna+q3AFjT3LnUdTAf/RyAmxkmOe2BL/dmrMpHcye5qYbdoNR82wfZySaQdyE6/c0mgi0KRT
WlmimNwZO+xmvR2x5prISuyjY2BYO/sgoqXwCT0A3/HqxOqYJH+MXWQYK9s6mDPIB9FzkoIaD1pl
g3per3Kg1VBkeEhvN20MuciEdfrk17j0UizxzjxtHgWarHKx5bpS+jKdyWEZON5jygh3NzTgUs8r
KJ9hHzldI0SmqPwgt8OE29C+zOWbnHDqwdkiAXQfW4RcLDSXbuRnQe6NiV1HLTMUlEVMaPz4h0U4
a1a4h+zfT6tGpfW+SibAVy4AANdOcTkIMroLp8Y8K4rxLq/kd+HFIS1Rg87rLUZy28JWTSgznVOu
3cx3SijB0K2/U4kwjA2pnAwheK0512+BzbTasKKS2tb1USpxdnCHvfTrClxy4cggCQK/w1kYGz0W
lAYMt3ySecT/3K6dCTuUjpx1T3hMYCZu0kNtCc13MTHhtFeFB3wlH2KZ7HJQm2MU7eySISOwk4My
ahPaiezOPp3jYaX5nEENEJFfDSgtotmfLXEqvqCvbL/WIFmJpsY76JgvQ11hkAkqbaUo9Zzldab3
X59lLQgpISs4UneoZmj8+h/LzRkZmSLlvqrfntd68+rasMMsOAcI1bgzHsGZ70b4AjgyPzx/aPY7
2piXnwplQbCaKq5cBcPbJEy6B8lMCktC98LKYRke56j3eZbh7RjIfrWXhzT9QUCUDBk3KiUHFh5G
gxkqBTkYt9erPRi+/BR2mG4YMmBy0tMeDG0BU7U+JdSfdTGrGuUdSt/BPDjZGBiP4QVWFWRf7BZ3
2JKp+JkbnNjPigU4uXa2VFxgSSYQDhSNAEM5ZQlQ80pezIreKSbnmsgsARvFVXQjQuHiYCuvYws3
VYV6+dWULWmpwmXCX7miC59XTlzgZoXRvq9jCsiCXutErcMCD9jNJL+4fuOQNG95vXMHB4sfNCv/
3iXFRnvEzGZAFYKuKySBYl1IUwiFymz844hZ6jgJIH4ucFNIXUx1q4gBpAHNSM6wdwtxJJAzYERR
+ncrFu/kCbPgCo0/OJ/XR+bIY9RYAl964YKvfh5t/7l2trEBlbcKYx6/S82NBXwtirZAfXqslreq
m05PX60bBtK9zPftRUnhyxWBk3KgbnJm/zEGnQUdcST698CTf6VkazXylpHeYUnV8Y3cvwBlaXe8
AKpavCWr1wiH0sBJ4Z9N0Bb7eIop457kBmglS9b7MDX1qbUp5NP6UORR2MR7R4qVmnDsKHo+GP17
PjS8DG/oZeVrBkAtEndio8EN4PVq3mrLY0ME5G0BzsBX1UySZMVFM4CGBbyxoxEEfud1p7jZz8ug
ceN8ODSQJQHx8KhNyHla4GGCImT79lTnGIDSKZBXPtDzeDA+5xS5Gjt9xEI+74NduT2cj/dmzljP
l08AiZ+RUYnSQmVbKM3XvbV35HScN47koYxEvOHxqCjjE1i6rkMhkqNKOVKjgVPb13jia+YQCb/f
AGCdpz9CtXpXkuWE0cPTlHT+petZbvNoqb5VZzMsIgs30DReK0ZQuEmD5JQoWOVZeZ5f52jznm4O
gjQ7w12Go8iUVfqzd5kQomKWmaQgw98PS+3GPGE3eYH8BSH+esHGh5ZJkv9alMkFuRiLdrFn7vmE
XHJf3J3GcEPRILarMVP34lbIJ2vAo1JBa4J/hP4PqQevUTUE9ZSRCs3HzEkOV9WiAniRgHGLuUc/
OEJI2zmsv5jFgY+6SZIuLhzSQDHmmMee0jPvRh7kBkb/A3d/FvK0gW5MLWogfHcDQ6hMKaTgLKAo
ymcFz7qD9JYc/6/DUtycer0GS4k8EWOlqKBgnx9NOCIZX5b4DTRf6ch0IqYuwdCnjZvl9M5dl/4j
02QP/Zx1AisMfdaKSB+9hhuR3etYAp+uX44h+23s5U2Vmi5zHJN26ZTX/npT7hBhrHX5fYWeufiC
46eDPFtgWxYcbZlKPk/5GMmfiGDiOJS6ay1P8Jyc9qdQ5EcjKoOGds5HNDiCYKcxwngB0rha1cw1
w71JTuZ8HjAFpL1LW7GN6ebMMefU1XQLdzD6bpupRQ3bqAfo7sheVi4ChfRhAQPz5kQl6LZ4tmr2
dEJpsnfljc3KSWsrUJ/J5LJSH4yg64EsfBAQ723CdyGVsabF0FK05g0RAeb2QTPIo7k9acu9FebZ
Bphc0qCtQU1aEATSrvFm10vB0JIXA0OtIzkDglEAqL0HbAk2A8no/77xRlBVlbe482I2YIVEX9gK
mFooKlxxoSzQeevPvACclUyHBbwOn8vG/jsEK3xpiVOpmczHQ0UPnVs43R49+ZJ3L08OwUGESZDs
ksi9Zpnf/ppvRsIcs19GTimgjdlr5tIo9evvF2RW+8ErBttO+xjJbQPlZU+3pppXLiF9fqfS6MxL
9mX/zT4wLYZ7TNbCcoIUmILuiXLod6arwDq1oAlN+xpygW6pG8YBMpLRB2DisRMJmeoC3Vts/1zE
k86+FKIFtZBhu67wXfyLR3VBjkDPA1L8G54SJRwmnQacLUuvXMWjf3TKUmaZ0AlnccV6G9ge5UYu
byatpksci8UOREnlnxBg2TsyxvZud6nQUMUxj8TxIgm1T5Ndss0i0TSy1XstFStbHogO+T+Enjuv
b9BklTV3vkaHGHOspGtLN2bdxQ5KSHKV6qNpvISCkZs6tOx/ywD/jRdpKPEDyhLvVYJ4xrj+zg3f
FVmfLXvgUu/iDAWFEH/0bXPQlDD1zB2dzXUSAzyyZwmrTAd2sgGo1UFgizTNcO6dOh+1uu7kKDIj
6a3gmq6ahahDtmdakaqduDbr+ePRpahH+5LnibCnqaaOG8m55IrcXEhU0H7qUQNBR16IThvxlKpv
v950FHQTfoX4+UaMbA4p3FiHRsSZe3R8sBFQ+6nF1usKEH7l7m/jscUIqVRpz5qrOq+KmOFB78Y5
g3+YALIvdwQApeEheZ6oQyaufFdVtYkDd1HYSZLm1QM5wOA0jzOSZ6OW1Hb5At/PfzeGWikBPK1o
qScA2N0Xd/Zui1opttgrvVzMoEUhhiTV9RWhJC9fiq3UJbjL25EwEunIEwiE600SQNv+Zkcdkkw7
M4/ZWCf5tuXcw0xCJARkHSy6uzaJKOr0y9kX2Ha7m+mgzVOmILLYHRVYVPOnjeYD0ih/3a6lLEeC
13iRkC+RnaUABMqtpjJwhK62dUiTLDVQbOozRAOhuXfZwN85ojts1B/MiuUmeFk5z9rjPFLZdGpz
2+g/ORTfNxwpwXLrsZsnwO3RqVmV4/461aSr6y7j6RttriSBqrboXUuHpASWxy4hVFY1jd3uZHRr
zmnwv3lJavvzIkW6Lj0/XwktUDIQHAUBm6CFKkW2ru177heC3HIb4fZdr9IASVY+0HWKHzBhFrrq
C16fMpWV6Mc/YN8VwqsmsNXB0M6cBNNDm/3RO7yOyxd1iBIVGB+mLwRqo8zOVDgUpMJMcz000rmf
kGqXadtT9HFhfX/gydR+9gVsacV8IJ1WZAwqFpNQMOUKfdyo2lYdz2WvYeNlLss3+AyzumGF26lx
+7qOWazoxssM24a+iJe6PpjNj7hvEzEEix+7oXDaZepsxXs5vRmJfjBIMUbuj2yrbXm8uz5BVQWa
QY57v0GDbUJX4wBfzZIZqbNm2Ym7eKovOw/onAdKY6rIbqYSQI7b8+6uDXyrb6alhs8CbhtL3gxR
nDvQ91lSrRscF9i9ACdOCsmSs8Z6nb6hkLCg7gK/ls1XrbqWr2aXInhYpRD/NIqfsRldHf87tw00
Xr8bOhHPtn6Kd+/sNtvWf9VH35mOTqSk++7vZIhnYLGIsWNnvpRGgEctIj50ph7YxHxAbJL9EzFd
c3k9dOO/vv5SDEmA0bpsUvSx6vGlC72Z4mLMqe3Li326newgydokqD9AQLnlX7zXFgddBX/lZejZ
jKrBn1o0V8VsKilf7bpyDF/kEn6Cv+p+IsYofrbBZMIybE/PVZJ7idEbFjsPpgoTwDyKeX26sqIF
qYyFsfKSSSGrr8RRP4wjKs2XsZikbRFMIV0kouosGxa+SEv+28N/GCpg4PFQDq/G1Eshn8qYcl+n
iRRbFmB6aVqq7WYK80SuP5MVucryulfKWVn6AoA3VPiz2fsZRGV6RyA13meHMnzn4v2AjWUcK0tK
L7vx/LfpkViNxaeGgco8q/7hOHPlfdF8KYL5fv8M
`protect end_protected
