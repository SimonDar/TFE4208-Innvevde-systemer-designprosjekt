��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8ez�L��C~�46Ǜ��b���l�|a��U~dr�I�nS�h�$:��;�K�7y��j`Sk���G+WEQ�p�X�%y"р,������	���<�]we��?��F��>6$k��m���,����� Pq� 8/�`#_�\�u¿�R1��Re0|����a�Jv<4���]���VhO?@�f+F���(�{�I��3U����o�Ū���x�:��-?�U���\aN�S����8No��Pk��J��S�OW���ZC)a4ܗ5.&�b�+�q�!lO���~6(��wR����H��V1�d?�\0һ����Z#���q�@L�a����%�,h.sΫ*;ک��A��*^k��K +��d�sf�:Ne��mD�\ ��'G]♸��̡Pɫ���ϱ$`�O��GY����2�PJ�)Ļ0�#�v�<��" ���1j�o�>ZE@�u�e�g��- ��a0j=Ny����v*��(
�&Z��X߄O�y���f�������I�����_m/Z�fQ�u�DK^�$cR6&�p�,;w��RtM��V̚��XN-�io�Rx+B|)��(��9`�;�L�}(���`��T�2�24c�\.�����@�(�V�%����z& �<��Z�r�Pw7y��1D�1����ډ��A�ºA���*$��i����M�l�'�&�T�r+"Q+�~�^�j!rqo�'Pl2�-�Q'��]5a���}�Z���ik�� �"��n��K��S�Nz47R�<����?���%`7=��)��L%�1�^{��޲���V������D���md���5��2o���q�AZ��e��۵"sm���L���JĝD�	Ɂ�,��woO; �{ �|����Iꤙ�bW⤖�=�^��&���}g�Q�!��ʕ��e3<z5}3��y[��/U��K`�X�ߘ�/�6e��
��]Z�U�o���2�O�l�?�W�'�c\�0����Yb)���w0}�~�gxyDYc+91,b��2DH����I���z��?��yNe$�u��V��!�0��Y�zժ�{�s��:yDVl1�k�.B����q� ��IGU,���.�����V��>#^$G,�Y��5(C�I�5��E�V?�� Ur����y \�����gL�Bآ5��ItD�^��B�M�S7ȷe���6�~��w�\']	���q)��Wޘ{z7z����!\3����ys��ҁ�<N�f3�����~ٮ�Y����Jԙ��U#�����q)i�9�\�p]��ݍ�'�t
��D�ظw��$��ڔ�`%9#҅uYۺ���11R}�@>��v2�6�7y�X�5I����>��Z^�]�����p������D�S%U/yW�ŚL�il��y���+xI�̓x��jҦw�_$�-�Oa����_V��^����N�Ykmц�8�V~rw�#��^�84��@hHV�.d�È� _5���b�B!a)��k�F�lj��f4�� ���1:t���̐R{�����`�u�*n��θ��P����GV{���K�¦�x�Y>�ݻNM�&~�<If!FY��Y��<��B�Υ����H$�nE�FǏ|����+����r��p�T3R���K�J�)�e����&x�f٣?r�L�Z�}3��F��������'����0`W�Ts`��v���7���J�2��a�WܦI�:�%�����q*��~/�^G���,�#�S��:ɋ�r^�S�N�˫u4��LZ�a�*�(P�Jg�5�	+�
����Ճ��yHZ�:�&R,�1ž�����邧��� �y/�%�JC�d�>�r�we�c���N6� �*J5�Җ�h�;Y����^�ߓAf`#�޵������NI�o��ǻ Ex��Y��Y����h�J�I"��ѳ��3���|�'mPö>\!A���{e�z\wY�)(�ƨ�ȅ��?�����7b:���`S^3n�̚��w1I����{�����v��hr!����<K�+�����	�M.�;��������O��YO[&[��mS7%[�Ę�o�j�TR����%�zn���$�8�߸���qsTG�ؘ�A��مW(�H�Q'�����*���d\���ҺU��hm���� ����H��GV������	��:t�<� Z�m��0J�!�DG�{!�➲L�<�L��[�*J{��8Z�9�B1�C>�N	�5SeU��n�0�M^$dg��^���MU�}T��(ֲr貓�ͥ4�|2=���H��[������C�h�^0��ؔ��-�-v��j�;�[ދ�z�O+g���E�L��%-��
�zB��x&�#���=�/��`m���	�g���HN��SP�C�(%������ڟ�"������W\`'x�㻕�
�.4GBs+]�Rd��{^{Z[�z=�V�>��24��ο���r~)y#S4�>}�Z�v�ƲT���H��wb1�)��H�c�K���Ng��M�M�r9�W�w��I�Z���9��}�.�#��%[.��I��.Mo-��j�o�үb�V� ޒ}�����֫z@7<S�Uf��3�p�B�cd��W�4^��{�%�eI^�r��0���ʖ[h���ng�X#�[:P�I�5&3x�iS��e��7��h[��?��8�5��Ǜ3��?K�͞S�Y�/<1�_D`l�z�?�:;IO���̪9�o��yD��P4�OZKTT޳W�5>Z?݆١�V�{����;��H����]1z0�`��M��q��b*�)����P���a�
��$ׯ�Yr1���aw9��R~ �G X];�~�`�0��rg+<�n�\�sOt�ڽ�ybڡԖ�ۜp{o�:���)U��촾@G�*D�!H�}ȼ�x|a%�W�Z�͛&��X�ޅ�s4�2"��%����y|1D��|���D�i�;b���X΃��^μE;˳4I��D(k��P(^��Gd5�����ē/����gA����Pw2�_:�n�F�^%Q[�^Z�4��$L����X�b�1qi��0��ݗ
��M�앥��������$��&���S9�w7Y5��\]�C�y��e�� �c"�J��/0>.,!�h��!���*�b?�=
�� �����T�������v?w֪��x��mU �	6��ډ��a�3��e�#,�H&q�=�R��j<�ٝs]6�Z�:Z���gk�1;���!��c�)9+�o!rυer� aAq��$*�!:��L�m�s�zF����=�G�c1w�e��l*.I�򨬆j։~�.y��k��q;uAȪ�ܜg�z�{�4����r��nא/�����e+`�K��5W&*e�w���%E�[���?,Ql�����+i/�V����Q�-��&�b�7�jQ4�6�Ev����S\�ƭ��c�'3/�+�O�C�o�,U�p�l�q�*�<4>�YPUD��S�����3��<6�t�+2B��ظyף�S,~��v��H�QmT%���i�u�!�'�G�G\;�����-��\�Z���	 ��Y벬�*[� �[I�UK���g��Pԑ0�J���p�ۨt��j^MW�Mʍ��f	���<�jw�҉���N��k�>�sup�+� �?�&�͇�owfĭhO�!b��)l�F�ٔӅ�ޚޱc;N�QF�&�W
�<��LϢ�����Ke|�5�Rx��?�]�{ŢO�'E	Mk&Hx���S�V"�!���vۻ��".�K�I����AE|`��S 9��,�R��X�	�{�OeH\��_����>��Q��/��h���ŀ�.k��\$x��oM�@��ږC�hFv!v�O��~�"���w�J����$$jbE���A�������3H�f��Xƨ���e�4���|)b�D;�YgGۚ�C|RGH��'��X����Σv��dq`�yQ����a��%������7�H�]�G\2�x_i�-Dve�/U8�&-P�*��������9% ����0��xRϬ�X�됪w�_�{i����]i�b�e���3ZZ0%����ǖ���}E2�V�Xi�e<���G��k����u����6i�Dqh����L����נ�������Rȃ�̙/���((B��/'�<hȈN�*-�b��ؓ���O��$��:D}"�K�yd�4np�&��9��3yˉ��؈�@V�]�S^�	�ϑ�:����*���A��۹�+r��O��ք��h�R�]��2/��dw`�-��}�^�i��W�?sP6r���e>�u���sh<��mZ,v�H�;;F�R�VN�����Ӵ�\@k��+�NQ��h�L>@P��l0̸Z���X,�?�~+��p������o=��;�H]So�_��Q�b���d��ݥ �+w2���!P�s���c�1���{���}�C�|�Z]M=E�M�����%,ER����աGɻ���e�撕�|�BdM��ZJ5�}����LvW�d?��5�G>��4�y��tF���\q6�;ރ�� �6-�Bڂ��5խ[�%#8#���0�u9��3P1B>��v0"l,�a���-G;�� �ԕa��_4�;�읛��V[��x�s�ND����ۊ]L4#�F�[d�mdz!�6�̈�֫�0đI��Q�tlU�}��sYO�΃֢z����`}N����,�";��oC�rH�<�E��V�LNO1��Tm��%�j�ep!���=-����E?��v;W���������JI���cj֣_"�L���{�Ԅ��گv��3.'�����xL���;t{��8;R9] @�n��<Ip��dl�E�)�b��#�.<�hx>�)�w�iD�y�-ǏմT,��Y*zr���dż���=����iX�G&�O�e^���Һ1B�⊐�xߎ���۷�U�<����W0-��GɅWa��3w-(\��{~_�BfS:����Z$�H��'��"�yv��hku��½� ���%A�ø�����c�"�#�_zP�5�]��)u�r���c>t7i��;��! �#m~/*G�g\��
��f_V�*@��(�����~��t{�������SK�+��]̑wv T-�O��v�#G���of��x��ک(k�σ�R	#7���Hx�
��ET�5������A����M�<�K��gGZ�D���ޜ�5zt,Ⲯ%F���*�-� x�a����(�,tm�y���RcSp,o4��A�pu�N���b+�l~Q �T�Tfz �]�Z������՘�_Z_C����n'�逡�2�:X�^��Z'M-�4즽l�6O��ʼ��H0fV�)9�O�	���J�ޒJ��D�z65�t^,��w�) ���^
z�ܴe�L��CٽEȑHí�=a��vw2��r�<�E�"��3[Bw���e�+dr���s�t_HYVie�A�X�b�nc��x��J9��j��˻+��������H`�����Eɲ�ӷ��S�b�.��(���PؔS���F�:����������Y����k�����m�Ψ#5\ѺOi8j^�fQ�J֙�Ve7�Aw��!��9�]SA�c�#*�8�p$0�1EK���KePwֳ���mҾ�%K��j-���,4�m��4�d"��s�c%���Q��<iߴ��k5�n,����H��ۑ���)7�S�.0
+��F�j� <+�*�T�I�FՀ7��d�im��#{�V��Х�y(z��X�}p�}�/M� �F�F���}�y�o^_+����x���Gh����#,�c��8k�ޓ[V���MV��u%��>�`��Nѧ���C2u��w�	_��9��N�dOwDݯY�v�T}�`	�2%��X�K��tB �V��� sy�����	�K`��������Y�]�2N�ĭt�wA5Ħp$�BP������lI[��;sOġ��>|��Y���.�)>Ԍ�:n�|�?��3' ��ݑ8j�ä����P�\�E�ӕ�]"��(&+d��dȶ��:�q;B�+]��˚���k������8ݭ�I�w�rѐ�ח�濫ȱ!@!�l�X ���6,�!�1��3�~&!GgC�)%�j�C@yӥ�;z���'Z�iIq$��0��GΘ���OF�6^�����o���˨ ������Q�)Wu.3_����U�Gɘ�ad6�@��I&�[���!f�Fqԓ�(9'�f��Db�d� q/�k�R	�A�Ro�w7�#���fVKVߖ��a$�9�\)&ܚ���4+��w��Fg�]\	�J<�M�ɪ�_P�}�~@��#Z�pVj�E|	"uW\#m���-|�~��0�tX�[����~5ϛ7�+o�ʹ8$9o��W�5{�&���ú���5~tM��<��W��]R�o59ә =���舫Td�u=�F����BlY�zP�h���o:�afĳ���%]����U�O���y��:5iJ��bޚfH���0��X���Ѫ�Ne�u�����^�t�$������WBe*H2�Ɠ���P����V�	�K���Jv��26u�D飋�6�3��ݘ�ċe|N#jc����%�)Өк�z/�"�������+m
�1X<���L��-�'�g)J|3e�i�w�1?J-�r���O[��eA��jd6�05�
�B��	���y7��~qU��d����w(u>�Հ�\�?B�<[%ѿv�z���|k��WFf)o�w��-d��}�C�5�d9�(�����gW����|7��(���0���]�w�����j�GґD�Hy�����a7��Å��]�A�hx���|d�8�_w/��Ie��e����k�� � K�v&�U�\��m�/Ux=���5S'�ުV%��(.PnI&��CV���f�x/�!ӷ�(q~U�����pz�4�5L�щ�S0�k� �_�H�t�ҥ���Lx���,@�K�h%�к��W0�SuU�� yMZ?��m.u+	�tf�<BMf>$�}Z�׌��,�@R �䩲��0��X����L*�Р,/���ŜH��S�/���G�Kd��|0y����=�ku>���4�Z�Y�z��y��7�(�A$��P�b��>X�n�Q45a^��8�`��M��{6��0��\E�5yވٖ�N�/�S����p����C��퍣��`rl�W$���<�9���H6h{r�]%�7W^�HW$W�.���:@�D�ݵ$���.U.X��:5��q�@�)�R������,wg[ �e�����j����f�>��|��Kq �ы�:�l/U���zrP���,�5.>o���$L��E`G��xzl��LfH���d��n�5���$8�9�%7w�z��/x@��U��;s����Y�����Q��Ⱦ�s�������,��$�LU���ѡɑ��U� %�
�u�u�ь�ࢲ_SV@S��u�+H��R��D����V�FGؖ�r�E|�)u�*���E��-��>��L&�i:l\o���b=�M� �wJU�W�bu:�y��j�A#�J�g���nޑ��jTfM|=)ɤTu�X��#p��������H�̿�l����)�\����?8I��( 2�dȶEr�q|�W�k«�`1�|i	b��t�=���v��2�x�&�Kp�?Q�=9|�CZw�j��e��@ƒ5�s>L��K�o��e�p�A���{QҰ�f� �8H�(K����@���?����"�iW� �G�t�h��G}rkY����]�b7q���mA$d�1�*"l�EqB�Kz^��Q��/V�{a�k����#��dֹ�;���*�z����ũ@x_Պe�`yd�:���M�}�]�}X��
]/���w��<=���N�W`�6�)#*S��<�	a�\�SPTB��ͣ_�g�НR�c4t�+��oE��ly@֤k(4>�����j;+1{�Ay�<��ΐ� N�X֞7�Z��gv��M�f:�!*$��8K<v�п�%�:Ь��I�p=<�x/`�u� �`$�����$-��ag(ON-�B�G8��HO`�9�4(*n{�1�a�i���6򬨀.b��a�s ��:ȩ�����9�Q��WA��H{mTA#�&.�|=���18��IxCM+c��.񢻭Ͼ���[D8��Hf���������Ś�¸�� ������c$�A�����<�W��=9�+�?j�߮��3�`-�OUR���@�1���T��cϰ���CIy��U_�=Kזj& �`e��l���2ظv�T��D2��Ջ�^�7&o��F�����&�ߒ?��j�n�%�~�g��B�؅�6���`O?�\À_��.Ѥ��>h��\�p��	�U�C��P�m�xQ���|��P$Z>O�	>��nhAS�x���NZv�Z:�*]&f��Z܆"�E��ѓ�Ut�_��f��"����^3�9�]�(��SE]����ИA*߁�<��Fy�i��I���P�Jp�����'�0S�2\b-q�{�z���މ�Z�0N���xn�+8�km
3�\>�3��Z����ZJ:`F�:����:H�m
򫓪pU�]��6{I�%̃���iCZÇr0j|�@tC��[�'�wGC�\�яԪ'�j�ot:3{Q�Avz[��"F�8�B�As���r�	R���g��U�@������"��/VոyIE'�?}���Rqvz��^_�*�6@��L[k{��|��c��Nd	�7�m�
%��\q`{�����lLJ-�~0z`ɒ��j��K�,��i~�2y�U�Y��&��}�����3K�l��~ʹ����Ʌ��ˢ��/C��c��^��v��q�Ց���$��<[ovw��۬�I�-���+��q!�E�N{"d�]�#�@F��0fR.�@���{:t��d�U�)�������f�	����{�MM�/U)	�AZ�B� Pe�Y��	�c�6O��D��HG܁���$����>�%��6c������.5:0䛎6�2�.��!-c)�~�<�D����dǂ�̇�t���9	 hؾN�o��+�U3��� ��[��;��HnL]F��	7?�ɶ}��`�@G��2�z�L�����X����H�1b75�tm��+��՚��BI$�U������������
d2{��c��/�m,�Yr��ܡ�2^��M62]W�:���n�x�ᄾ��o)WOT�K�Y���C�y'
�ɱ�V΀�}����He%@�h5�ω ;,���|��kq*&6%��Hx}�]Z����ea���y�P��E3��4���F	lX��0;v���%�.�0X�<�C	��#B) �G���L�j�
���#��"�[��o�|�P1�
�h ]��Q"�t�K����W��/s�L�L'��4����GJ�<��z��O��!T����=�%�}֨{�#�´��x�[�o��vޮ�^),"]}P7$=��C����̘�{��zF5�AO��qɸ:�������.i���8�Vv�?FPt8N�>�^/� \Ns�ǿ�(}є�w��#]��sbp�:g�5����X�*@:���`�3�gi���q�ܱA? ���ິjP	[��v�]*�a%�#���J�5g���H�
�Jt7���C�O271�����>�,��ze�����69��["Po����k��u3{�(�7|��]�,0-�Z��̱a�Z�>�[(J�>��g�c���VI��5��R�Q���t���^=7 ���Wc�Һ0Ղ�F�Nh"87u'pi`������-^���Z�Pz��VLE�ۑT�_9�?1`Q�_���B�����k`;��6V�����abqimW�&}`8C+\�#:c��S�}$ds��̤�rfmoY�	|h!�|���3��7�4&���"����LO��V!���|����%U\��y�i�A�fY�u��m���c��^u	���V*�t�}E��$���lFݛX�;�2�=1S�'�*���9qsg��>�����Q���h��5v�:Ցl	�����c� a]M%���/�@�:ڸ���,K3n|��l��0���>խ&�]��� ������!`��A�댸���g��{����Gc {R}vtv�*WX�j)��\�:K#̳;.OjU}8��4{F������r��qpl�������Y�9��L��g��A2L�^P}'-��Q� �e�Y5�x���M�rw���}��9�vDqˇ�&��
&���}|�wP3��7������C�\����ʔ���m�����T^�KSb0��T�X.ڱ����=te���V-hvR;h��h��%z�30�Ǵ��_�F�=0�|/���쾺��-n�^���Y�ľAg/���5��h?+�3��q6�YO��P�q���6i=�������]�WV�L7Ğ�����P�{�S�i�["�{��o����xi�K�z�^Ը[�BF���i'4�%H�5�$y��@~V��z6���j�-c�m_���n�d������}�AH�<����dp���/B�&��;sh!�a���_�wO�����Ƌ&\&�-�U|@H��g3K���0M�#h���}�K�,�x>�8q����'�@�H3�/-%);@�&��d�����>����2��#^�����v���8���#O���P������*P`�t��2�П4�S�D�8��{>f��2Il�a�t0�5������i\�lY
fq/loh���S�Ė�����b;y�]���i�Ԏ�S\�/Ձ:;{�����dǡC9P@R�?]�X�#��;`W|V!�5փ�#ěe��Ɲ;n�:�����=ރoe@�K�H�u|��ȕ���6�P���ZG�*�V���O�4�lkBѰ�Vb������,�ѥꙧx۲Đ����w
�@�������T�SWf���c�]��'AW�	1�����x��~��uZ��v��X����/@�.���=y�OR採JX]�`Yo�m�ե�^�������Q/� ��Ӗ�e>�FƐJ�����&*�`qު�?�:3Z�f�b���uh�6?Z#�0+��F�R�:5J���-}j]Z�+w���&��o6 �[N�qk�H#�=�Oarea�E0������N*��ܳ9��
�{��������n�<�O�̓�g�ܵ�)��c��ݡ�a��24���Ų�p'J��53
*<����8�k��af����;c'�r&�w�v	M mD���MW�7œZ'aM�\�[Ę����S���A�w�o�Ms��܈� ��W-��!�E�u[�[�x����z2��S����Y�2����l)����_ҿ�j����?^	�����=�8 a��%ړ�8Ll6��=2��U�TJ�"��Dni÷^���������SV�MA����ߖ����q���}E�����P�ؒwB��$6���d"����'�6�ܹYt%Z��wy�\����k�S�D���A|a���(��Z0'xȎ6ˠ8]eZ���SW��A�7��-[���	4�T�1(�9Q*F�vUE[��c��6贤�0�n3y`
R�6VZb_�V�=v�^z�&�0��`w�S��EB�؇!�&�H�$�&����;5��d��~q8�H�ë�_�BhK��z2_�b���z���46�oY�!�a4��QH�7�tfx!U�i�9���*8�UY��h��oD\47.ϐǨK��v�a�R��F֟2�(�t�G�{�Sě����Iy�B]h~ߺ����
��P3{����x�L�a���!���<���o�ڳ��
W#6���V�L B�u��q�Vh��Zw��˘f�������n��]�&*�F$z��,'�l��UaW���I8�Si;q$@��7�ƻ���/՝�*0<o}����>~�r�����eWx�-$J��Γ�P�m����P�Y�6.���B�~���k���Mr�aX�v��h1>pj�'@���џ�oK��ʳ����}��o�Z.|�eKW|�F,:��/��Ȑ����i�F�>w�\���Qy:G�����>�u�7b.a��1LϷ�t��>�oHƕ�MX�ŎG���-�m��E_�o�-���,s�H^ �**��$�%��A�(��F���l��c���5�������+I� �A�,A7�wP&&�t��(��.`���3�k�L������X��=��la����3�6�J:˫9�pt��(d���
�9�D �ǖ�*37[���U�����A9T��^�k7�4��`��}QHK���ӫ���G��?���V�s�X���?��mh�_[\�ᴽ���<�ݼUuch,�ZZ�jDC�fd�B��n��d�:�da'�9�6��mYci�M�V�X�����Ki��g��LgKi�<Y�&���f�G]���N��g�4��b����:�^J9�����rz��P� ;������{ʔ��ܹ~���hVkj�F�Õ��ӓ��/��Yb�X\(f���&�����	�G�������v���F
��o����>�4σ:���/q�����<)s��Q��� �j��Q�,vn��JU��F}U/U �zE蚼Tm��pSR[㾪�/w鹈2�>���ȏ+�<h�狕�~^��#8�i���b�8(P�U��g���u_�!��z�Q�����G8^�F*6�S�Ы:<����xol�{�G���6D��~-�'`	?\t#u�MtC��βLB��tW�J&8g~�u�3Pk�xn�=ф� <��@�fpnƼ��~FsU�4o��,E�/�򜷟jj�&\�$-�,�?�m�ӌ�6�/�UȲ!,���0�(�P���FP���p��'��7Sݫ��םt5�(��]
�(n�Q�2�7�yY�b	����]�@�1�o�8��A��k��^����g���h6�Dc���9��z�#�n-�i��D��b�"��F�"��N��|���$r�w����iK2��bQ���=�#c���яHO�⣀c��e������l��r�8����:���j�G��5[�m�8���;��ڬ�oI��
�����;�����t�y��J�Z4�x�I���p߻"=���ĭU�kS��gA)�xݧ��mXǲq��&�e�����
NO\�RS�H����e�xc�3(��$ӓ7F��TJن\���%CV���s�D�Ʃs�.<����>}H�A]$�'@������J/��-�h�z�sKɠ.Ԝ����%'�s��C��BX��`�F��	��W[�m`���)�nj��̎�u3��8K����T2�~�=�g�xb�u?}Z8�����-�f댖���&dT��m�r�\�崦�ȏ������=�����i7hρ�Bw���@�2���J/i<Miǈ������JtW+`����[�L�׈�1��v�׬N�*m�Ӡ����rC&��C�����K�p0,nZk��Y���k�1��{��E�i)&l>��|K��X]���8�G�r��y�W���@x��a�D�ʭ���^$,����7s�����e$S�$(�f��#ۗ�3#W��/��νc���}�/D3q��FU*�#ٗ�i��A=��Ű��5c��{��p՚��`��������\f�V+#A14q��}3�� R�CW����i.@�5{ӰH4>Q;Q��D����Pc:�7е�=�Fq�Y�������<Ka�J��\|w�ƇG7s�|�^��2|C�?��7Z�
���@w|K����"/�J?�d8lz�� u�A&ȓwk�]e��:W~0�&�
E����V0D4���$�CL�t��nV#�S��xGb��z͌�6	'\#�|4퐦^zvu���ܑ�RO�T��\��dj̵r)��=��ϥ�^3�����le��NT�|P;��F���yޜ��&ܚ�GVc�w��=���D w��Rp3x����̸�'�� �(����H������E�ߑ���	�F�0��6��Pσ+>FA�z��Ӄ ����,W
�,W$.�c�j���� �t-��t0�����PK��P��|J�>��	rP�}�t	��H$��+"}@��r��Ɔ�;h�K����;���2�'��7p���w�Y���j�~`�?�I�w�.q��Mb���t>z��i�ч�(���@���%G���]��_�(��ĵ��
2P�r��ѣ�z�۵#�~�
V�*�D��T;f��g��4�sZ	%=�����|F�0��4fX���c�XH��u��_��	��a$�$��\X�+�d�W���;`�{�I�n���@��eN^��h������:��)�E�����I
�Q3h����9Vy��l�J�H#��ۛ�PgC��,��V �Y�aNb�%�?�h�'JS�9I�n����\�8D��V��_�7:(����t�;{���{wT���c���/��_�)��vZ�'�{<e�t8/{�G���:�@2b�<b��
)�-��m�t3�a�|�qv��L�pk��MX���4s��Y.>�ׯqRBr��q�zZ�|ʬ��@џIQ�:�1�S��v	�+��I�#��2 v�+T�g;&gt{'��
����LPC~V[��L�'^!�J"�f��`_�Z���Z{� ͌��f�#�$��C����|]B�\�e�Iӕ�v�a��䋢75�5�m$+��OfBPOMgԽ�!JhB.5>c�:(�R��]:����8�#.6�{lB�w��F��y������en�_	|�os��d���Q��R|���@U�!�K7wM���x2~u����Q4G����vcj¸�1{��Fi��	)|�P�'8�_�?]�Ċqi�%�v|m_/S^��u3L��r�3�C"��������N��pc��ϐ����"��-w5	D�Q�U�t�}�9:-�����`�P�S�:6��4�%��)��c��' !�D8�	Y�KF�i~ӂ�i���J����)da5Ccz��c�E�R�-��dQ���҆�R������E�C��Ё�#Loȑ�ë��@��~W׶N}�������W�p.��"��ͺ�7\����c��у����B"ÿ�ŽJ=��ⶱf���1N�E$�c�8U~�U P<h9hUE���A�.�D����|&/'�#y���9�NP<&̬�D���6� g\}�0A�<�� �=�	� ��ƭ�/�z�bav;�<�-�4�̀�h]ݟ�������A�Z�-��	������%	��f=��h�x��f��`D�X!��N6�"?Wª��3�,HK:���>�l��m�ƶV���1�����#��:�_r��:�_Q��Y_�z�6dH�A�J����D�"���F�C�#������TF��9�|����~��%s>=�c&V,�2�����]�G����S�
P����|�T��L.��C�ܣ��&�A��IpPu=��]��Xzq�) ��B/��h�u魔/�6���E@��� ����晃��p���7+p'4o��d`�ԡР�����p�
#_����O���W���:���uw&x��ؽ;�$~��l?��kwfQ��kA��Cv��I���r��y
9�r' �erI$�J�X��l:0f��*s8����2�Y@������[��AS��
d�ސ>�]<�h�����/���a;ub��������
FbA��Wc��A�*�c�X���h(X ��½��2!f�N�7�M5����oG�jRF��=��-͑���O��+�(�:WI�w�t��@�h��^=�@IV�ĕ-G��v V�p�����&{���{�y��#1����W�N:F����S�Z�9l����'��Ք$Ѹ<Y=v0w�����4�w�����ݻ>e�.�|���Ѡ��j�-ș���S�b��h�MAdˬ:�R�#)����ΎF,��	L��e^�E�f�"���8mĀo2C,���@�
�tZ�
�[�����O�φ2պ���[-EHqVXe�\ηмߛ^�^��
��Q��҇&��6�Ƞ�H��WG��,�p�"�lod�r:��$��ς[��MEi�Y4���)=Z#Y��(�;N��qY��K��f�A��!��h��V�dNv����2���`<%��6���D��2,�N���܏�o%0r��WA�0��M�&���;�r�FG'�b�~S9��j�F���m�C@l: �W��q��b/���t������H�)N<D&b�B#� �]���V������׀�p)��s�T~�b�mՒ(�d�'%��N_pV����g���z	v"�,�D�c����?y��Y|[��'���r�5y�ts��>�͗&�h|��q-��ԤM�Pl��`�B'��(և��8�｟z�o�{�C�X�kx y����N��� ��SL��?g٭��n�/�=�,l.����^������w��p�Fk$g	&��I������(��۟��i5\ ^lh�_��%�gs{���G���͛tY4@(}���棹W�\.J[���g�e7�s��a#
$�(��ŔBB�0k��U���)KPJ#�_���ꍃ�=	�"%����]���/�`S�;�@�>����)��d]�*�C_��n���RǾ��j7�d
+%M�h���#s�Y'Q]���;
�~UU��3&� �}�o�,���@X~0�=*�Na��P��UYw�W�"r��+S�4���Z/�ٙ�\���AB��0 p���'fR�K�wy��i@*Q���'�����,I�Y���~�')���Z�3Bt}���!��+����]B�Ǿ7�w�bvn�py���o�{�hk���|,|�hȓ�������MB�bh6W(�	�>dγ�,�%0�=�~��&�
��'���0�Ct���(���f�U��o����p�i ��U�Oi&��>k[�t�V��t�"���(��`�|�s�:��jKB�ݞ��@yͷ��ju�*V�T+ɾ��W��7!{_�P(1nV���H�s/�I���/�d�����p�����t�$��#s�0�w!DGd	�}s�Pņ\�ڕ{�@4�-w'��3��Í��z���jYv!#$�Bt!��X����XL�����T����SLf1�n��D�5�$� �;A�/�6;�kb��%9	��Ǻ~\��`��V�dRk�pUD��+jgw��2y /X�����q�����Ȓv�����A3���.Ґg�J�#S�*d6-K��Ժ����h��C�{
�Y�-�Ї
��� �C�(��\�z7��3�o�oA/������&#/_ǳ��3w��ඊ*|�o@3fNٓ�"�Qq�E��*��U	�w ���m��2�����̷����_�p,�c��&#�~P�[ҭ�<��!kL�2��Hzp�96i��Խ��E)�;\��J��/��{�`R�o/�$tUSlX�Wl�<(S�Z��݁���)��)�l�)����`h�ҫ�1L�bqo�R7|'��?��[�K��#-��b���)ƿ_�J�����.;=hq�oFX�UL9�ˍ�A��0��OY��#�ȵK�Z�>u5�Hd=\�<�,����3|�_������#���dG����ȯ%v!����]�Ӓ1-�8�"	�.��`zN��ʞ/j�NB<mo��g�E��s=9�D[��B��v#~Y��!M�]�_i�PP3�lY�4xĉ�uWf?-* /ła�ȧ��i+��������ZH�:8�c��ѵ��Z�!�
l©6�v���,�-�]�RF���y�K�cI2��gCX7���j����
U8}���&@vozL�E4_Z��B˷��1}bjj�q�ĕ�?�1 TS@&���Ǧ(����7����z�L�//$A��"�Wg`,]f�U@���V�a���*zP\R��*��XV�a'T>Y��!:i����墴Sh�L�ځ�����v^��O
�r��{7�Z/�Ş�{yK�ώ��<bi6$�� ����V�1�|��a|*r?�:����rxD'�Lrd�<�	�&l�Y��Wg��������t�uDR�p�	k�}�|{�=�)�cF��yd�D�F׃OĪ�/ak-�n%��+�5��o?�S*��j���@�:=(q�<B΄>(z!��ב������>�#cǃOT%�7\�~����!D���5��b!<����230��x���@��]L?69�<X"ȴ�;�9� ͵Ik�]t���$*Q0����Z�rrc߾ �m���O΢����7�3�2�@���9��zm���!T+��,!�������t��|�Wxhqx�-E'.�ЭUU�xy�֚��W�C�bW��?<[%x[-��.��Cl܁%w����Ѳ�Ң8�����T�զ(��������� *���/'���i�:zj)���$�;������T���};�ݻ�<Q�Q@Ԣ���U\�Q�y��H�Q9k�XS|}���*Ͽ�뉪�Y����?���n�	>�
�M[�&��\Q�]�Y�+	ξ|�^�89��YNk����#+��e���G^���[��Y+�5:�	|�0@9Hz�y�+������t_������1]|�v��J�2ed�v�T*B������f�mT �o=��t��y�=i��D���U�"^ �xY�����C �ޛ�.G!������_��a��h�\ԏz��Gu܄J�z4XB���e�	��}>�T�W	����}�vy�U;�	i*$�h�f� Z�qǤ��\�=�t�;]d�����R2P]>���C�h��zx 6���FZ3���CS^xC[�El� _&brׇ���9;C�\s��T�Si�C|2_B�1�}$�:��
�]�ھ�p��_*��ˋ���y���=X�����k�7�@����خ�)�l�
���C��Lm� �@���1� v��Wi��-ȴ�����"��>B���wŻ�����K~k��A��pF�c/]o��_?��ߩz/xTN�v��6�;���z���IE"�k�7?�(ߍ�w2�j ��Y2���7�`��c��N؂!VV���U&z�Y%�(����� �2_�8����h=]�ò��?��b�\Ƣr�Pj��3�CLE+�v��+�d��Kߘ$��&u6�6�uN��0:jmv�oOB3X��+�����=Gk���+�ĨoE�y��`��:�?�$>|KVG�}�K� �/l֙&M��CA�_�����M_$*qqX~7q�ˊzGe��f
�ǕG�K������C]ہg�w��Pt�(�W�(�\ioya�߂�Qa	G;"P$�3IB|~F�Pn����:?��%�z�e����������f��ZQ�4h�L�d]׌P:�$)��pZTMR}j��.Ց)m ��R���I�"eźH�+��y"�M���7O�'���X�t�E�/�ĭF\�0"��>������HH�i��V�Լc$��t�_P�锈���
u?@v��-gCR��B`GXU~�� ��+�TN[����掉���ˤ��j$�AؙY�3�����<��Uk��TQU"?a]�����?�_sY�B2X�z.�=�Up���ty/
,�b%=�sn��q"�
���ha��_�AձQ�f�����U //M��F:W��C#��Ci>EPj��j�\���nXiC��˱R�ς	p�'�Fe::�i� ���5�/����2��d�ck��F�%�����W���G5�(A &w����#�n�;�{ʒ>;�+)?�Z���� �0������3i w�Lքr��(�\�+2��>Gv='�	�����Z��Vt��ʃ������y]��%O8(}�y!]&/K_kN`��i��hfc��h�e.��P2qM%��S�Tq��"�����a���m�X����K�?F�W���P�I�?�]b���%_�ZE�]�.�XAj�F�8�*�=-�1!s�uv݅Z��#=j��ζ������6��&fc<�hm�i.�P�cgM �m�����J��VlY�i��6`'�I�`2����q��t��=%�
7�"�^�L�,�32�����;А�(i��Ne�.v�ο�������A��*������t�%8�e����E�[�_{�E<HKC�@���U�m�^�ձ�+ey2X���p�*ɏ�󛍕�aC7L_Ú]�[0c{\'���H/���.<�xHzƾ{�Ǡ�H⧕�g~QL곐.4��g)O.}����9�*���o��� ��A~./5���窮&'�>z�b"n��0�
T1A/���am�G�G���W�G=w��;�r���US���:�׏���+�q�R�p@v|�����p���b��FX��\�N~�(�����9���h�fYi�����C1fPTT`�f�/���p�5��@�b_�_���V�� i.ּ��S��i�L�I���7�-hs��g��f�=]Z�rۥ6S��U�����w8�Bvc�(��ݼ�DX�p�˨��Q��J�񩁣$���,�	���124��*�Ja��cS�>��_E�Ot�~�Kn4l&ܡN�TA�HF}YD�~Z�>���4���O����*c�0�)��k�?�k���2�^��ɒw���������-�l�.ތb�G�����S i�%��>_��h�\yq�k��Ci܊�B�1�?(eq Ǘ X���r!�$y�Q�m?���۶�3,�'��	��?-�Rk,nx�yy���+�o��ue��O��( mꂬ0P�~��vt�ª�$fEV��'ot�ܾ�C!��M�䂥}N��yGi��e��i'���=�&�v&%��M�`,��Ua�F������Rzڱը�qq�F�PKU�:�*��ͫ����(4�ԅ�֢�����@�0�J�c.�0��5Z����A,%��3t'�u:�߹jX�_��ϗ@d�l���|���{l�nћ�D�d:޻;�`�@{v]�5�D���x��+�,���r���� �}N�&�;~]�4]���[�F?`	l��uW��[�a�ς/Z�݉�.pP��\C�*�s�깡8�UW�<p�G���F�����$j� Bjw �$S�5J�gL�k�����B5���hz����w�NP�J�+��m���Ҋ�^�!�l=�[O����2��w�G�k��?Y������2�[|�vOBce�,Z1 &1q)	,�[��Ѣ�����<��uS{�	�ӧ�m���C�Qxχ����o�ׇ\4��dh �xCd�21
��vP�.�F�rF�ÆS�� �M"J����\�o��%��{d���	J��E��bb�.r���K�dNoG,K&�~�=��d�+h�a��mgh�}}~4AhJ\9�b|O�o�'�tl��[���Ѻ�$�M�	N�3��0�1Z��r?|3隶�@���c���Z�Ņ�YC�g�U�UZ
K�0AJF����GHr��ADQu����>z�k���q���dj�B�G�!�qC����
���{�Ȭgp��Zq�쳅�6=���W7�}t����
��0;��%��v�:X?7�!����w���;�����X��6ÈX"�;Y	��1�$��RZX���)Un?������nN���D��������P�	u��W�vF�:J�u���>gr ��Jc��q�m,�Ek���m��q��߻O�rT��'��Q�e쐔�5yذI�<H�JyeJ
��+��R�����t���j%�eF�4C��7Z��y���ɴ���� ��Rn񗗙��<����BC<������ao��^�r>�R?Ur}������4��Z�i��b����,�Ed���+�c������k~��|�<b'�AAJeLA�����V�d���]L�j$�*�MoX��	��X��|Ii��Z2��g�h�lF��ƍ[R�o�����e��*>�ĩC��N�p�>�拏��������	T&~�Г(��C��;����D��"��Z](͕���P���,�I��Ս�9��(��a^�{�^���sЉ�р���^�P���&/���Ѣ�*���Rk!ʝ�������\ws��k��
`ʊ�_	h
��cH�>,W�1��:���1���Ҫ9tU1�"���f����"�Ae��A���
���=K�|�V��ef��V'�/|;@�����0������i�P�-7�P����6S$b��H�$�n�t�]��>�ֺX��6��=�Q��毲�|:.�l��FY���B����������Žp�ibo'S�t�eU����ۋ�04b����$�� ��T����g�	#��"��8�T3\��U�����u3�)��!�}M��ݰw�9���.\Ӯ�E.DL���1F3Ṭs9�<���i�d�^������S�s��ͬ*�2�9d�,0W���9��@��̈́©B�8��^�Keh���k�T��
�5w�i�+bY�L4���#��@\=.?���V'V�␤�C�c�.c���<6*�Ê����T�����j~�� "�m�� ��U )�<������0 �����|:1?|����k	]�حS���=�*��|�[�V�ߤ"�3�����T�,Q�O�r	4����M`�|�~�P�{V<�fI�:��/9�Ъ����������NʾNKx2˱�D{�94Z\��1j,�@+z�O���??��3�҂18�[�Ϳ����1u9Ś�,�@�%��c@����x�]�Y����/���r1 :RV�'��
���h�\oMR��s1��O�;h/�Qj�F�x��e��5��	Q+�n�)^�w�ۛq}w񸁓w��
�q�"^6+_?��㚕D�U��] ��MDQݳ|٤)��5?((��I�f�*�Ik�1j��\�j�l��h�褯%*]YAk�\kb��o|��^3�؆�uy6���X�7�U�W]]7�y���'�7Na���O��9�� {s��W�]VZxR��}s�����������D���GKlmF/>����Azn�t��<o�`��T9K�~�;͈{E�î#N��[#��� N>����S��{��e-����b�ԍeT&�/�*�,jG���Ԍ���̴��(�P'g��X�
>B��%���FbgT�A��$��� �%�B���	ޕw��@N�-	� �  ���,3Dl������T,������*���Se���;BzF�����d�PQ)?#�0|�}��B�Q��0a��u�\����)�&|E��k�Z����[#��9)��]B��tI�<�mb��٨V�M9)�5Z@뿶�ְ5�S6�.�f$����(O�����]�� m�h�V��ζ(dA("�5����~��<�b�j0V	�F����,
+m��|����v��Z~�ڂK�v�G$��u����h�-�?5�����JƸ��r�4l'q7��O�1�k�N���ߖ}
[Q���G�����W�Ӆ��������s�u��R_���n�'
ԒJ�YT qD̼aY����B3o�K&�3�m�e�G�`U_��&�-�c}c�[�TJ!'�����wø��)\�Έ�n6��'{WY�a�� �*�r�Y��7���
�V_����ݧs5K(G����G���Aݙ�=aG#�ڷ(P���bu��]�V#���A�����!��\m�b�N"?�sTbӠ���}��8H�dQ��b&��������~��d� �3�K�̘Z�((���.��&i޽I��-�#�4V75%	�����o�'x��H���rP�mw%�m��`�*?>K�/4����<�K\��v=X���kU�1m��i"~w&�Ŝ��[�Z�W�P�C��-x跿�V��M���%���4����/��>�|��5��#? ��q`��P�O����ĸSY;Ue64\�^��Ҫ#�,69�o#%lv��Qm�G؀��*��Ğo����KN+e��&)P�!��D�)D�/g��Jz�,������0��(comg����Ʀ�^��qo�n4�sY	��ڠ5+�9�Թ����ߟDw��Čﺒ{�Y���i��@ˌt�}�<�6g�N��<x�y�I-�q��0h�4��6�`8/^]��IZ��Ȅq �����ddd�S�@�Z�rGip�"YR���x�<������Q=@�o�H����_�H����rJ!�6�B�Ana�d\�4^��B���p5�@�&0��D��cʒ,��B���A��l�1�xs΂�*)@�ju��pr�Vb�A����:��ўOR\���q[�[������ �Y�:	�ԙ4~�%9�ځ�|�ȿ� W��3=0gE��&أa�Ml���F���+��7�U_���m)�1�H�#�͆�0�U
�ު��%r
uDH���w�͸Z���ѫY.Ӄ^�2N&�ƕ2�v�C�T��I��y�PS4�� ��*���ⶃ~��'��m��,�ntN��m��ou5�3�}6 �D�=m�]�(�A��͵�N_s`Qőb��̮^u��?�������8�F������M�#H�����Q�<�I��0^շ�S�J��K"��LS��C�4;��3*<P� ���&�׉��mVu�����(ۤ�#�+PS�1;Lig�j6H�$�S�\+�""��gn���p�J?�d�)6YD�t�v����1]�"�x�]�w����ݶC�L�����C0'T(5�x9�"����A�ϯi�L9� �[��A�"�bA�C�a��x8���Կ{O�0M0;�[x�{�W�s5��V�����c�EҖh��t�!d�����AX#\�ّ+ y�o�<$�䅲�����J�s/ʄ��;�1=w��W)W~KK�ҿ�� +�]�&�GOe�� ՘S��UI������eq�֯ɋ"|M̐�j�K���6=+�v�z�*�;&�� ���!"2:#��o�0���뜁��0��R�O9B���jvN�}k��o�}�T�xk�Y�C[�ѻ��1�Z��O�D;b�zd3�z��,R|�0V�|U�)���xܷ�����ѽ=�ɰo���ZB���V��E�ݘ��ϱ�NZ�ܐt� >���?��i�ܸ2����o[���~�Y�	3W���MJ�E���eur$MHu۳�	Q�65G\����w�:��#����h;��i��{�vtw��}�eG"�%?���NF0�!��W�yK�.�<œ��tmg�$���>�Bz�_n��Gc�/�3��k%����x��z��0G�2�hU�m2m+�����W*�p `��ʍG��$�S#A)�a-�d�\|T���W�4 +x��$ع��]�Ư��Y{h���Pز	�DgH
0bg����wVTD�����[�4��Rg�v2޿�w�
�S_d�'���"�u[���Ĩ>����F�	׺zBi��ey���U�C�S�"��](�ϝR���o��xY%����yC��-=��ߚ^��)���T/��\�RT��!ul�C��8E_O�Q��{"�d ��f���F�#�;�D���)�G�I�/� |Z��|�Cb���Qz����)�J{�VF4�kd��S��>�}�g��b���	J|�H�2�6I�H�����+��ڒR
-e���,��C�J:(u0#��!؍|���L�ԧ��3AR?6q��B���1��x�� �������:�ӦB����+��w����Yr�6�y�3��?�@c��n�r���7���#�k��<9��b�*�W�s�>�\��y_$�D;�gE���l��^ٿ&�k]ε�����!�7Oqި��ͬ�0���oAFޠT�?蜲��)-�.�W�O`a�;��ʗG �x����'_a)o�O���fcly]�yc����7�q}���[�8z�{E�cE8 �tݖ��C7�`^7{��h�h�*R{���8 *�S�"{>A <а-�N+4[k�9$T�P�����98��"�B�oV���Ē7[��� -21ʪj��K����b�C��pa�[Zz/Ww�)3��J2����l#��5:縰���4���|I.<��UeT��0yTO��܏��<_a&@I?ɤ�]�۽�`����+���v6L���8,)r��k�4 ^_3|��1Z��&]�',9��lK�x"�j� 4�.�ͽ��L��:~mr'��g+S�C����eq�`�S.3�S5ץۯwEߏ[p	�E`��?�a����	X\��n�`�ngj�)�{E�Rg��_D���~�ȯ�Z��mR�T��J�;le��K�
!S��U�m��]�T�M� ���KW%Rh�@Q�ɧ�񋴘a���$�l�9�ߓ)G�_�u?"Ju_�� w
)�������=��g>e�5#� B:u�ト=G�ɹtqm����?u$�A����f����^��>���<"�de�T���\ɔ�����)
����;ٍ�K�]�,j�0�®�6���]~���4��n;Y�ǒ�Et������x�}���{�h�f���t��ѽ;$e)��`7�^�4`C(y�[���τ�Z�г�0K�ҭ�PR��d�9�y��0��f�M�\(��@��C|�M�|@�ntj�r ����gm�;�G��d��7YK*̲����02a�� @��"����	�0�
4ſ7�R�2���xS�qRwn�To� �ʑݨ9I��NT�������%9l���/��3������(�=F:���1��=I�X �%:����G'[|_'���^�(j�^���oG!�9m�7��p�>i�̗��aM��+��A;�V� �!F�����e�W�֥�d��B�_���L���6�6��K�	��ư��,Y� m�m7^���QN�78��8~3S�7��O�Ӫ!0)@�gk���������߁0 _B�N�d���5X�>نB�`w��Ȝ��"�|�T��Ô%'H?�N%TF���ף�x���8�� ���
��A��F�NCWK�~��,�hO�|�d�{������R����*����tR�(bk&��>��WҞ�����:������V�L�S��yՏ�pG�~X��v�R3�E��zH9O��-�0)�⟱qa��X�������,􅼵��U�?�ծ�&�>��r������h��]��b�m(/=�QxET�&[N����//�c��\5d���4z5�v�~�ڋ	�a���3��	<�i����Б�!{_u��-i8�H�(�Wl%�:	�V�Z<��gߧWg~ T�+K��o]�I��f�(�5"�?�	X��2W&!t�w��������Z��_Df�x��hT��1*���T�O!TyqڿI�{h�jp��TcVTJ۪��%����PYjoa�`.L�4=��gMz����7?��*؝c�,}}��V������ޗ����W"n���y�M�91����N.�4�b��D�lV��3/󫿏+��H�htCMN��n�w�����JS6|���*� �q{���g7z�����U�E��)GΣn�3Ǩ7�sr� ���� Ͷ�j���!?4vj[��/�dߘ?���EgT�l��צ�W�s����XI���k���'�I0�"�	��f�$N��^����8�K0
v(s������-��na��9ɞ?�3d�Q�פc:�a%ي�ԗ>ULm�خBB���ޝY��.e|�WH��4�_m4�_S�����{�[�?D�0.��4]��e�6'pET)�[R;�2��d���U$����v�ڕ���l��8�+^��-+��7Rj����/��	hn5K5��O]O?}�÷�Vt�Y���Vg`wr�U�X��2�f��f��e�-K|���*区l��W	s�����.�
�*�$�r�OӉpf���g�a��R <�M�f��l7�x��(���3�|&qrЬ�9�뢖�� 2P�g�ElT�^.da��k��'��'�NE�'OV?ʱ�y�v&%8��׾˞�oh�Wz��~�?4�"�������"���7cI�痊�sɼ-�s�B��JM��o�f��œƁ�~w���S�ͦ��W�2�5v՛3����x��"��Q2������r�V%��G��9�.;������c`�#��=�Wͳn�N��j^��i@��o���B��,��2�ž�z��选�23J2�)���$X�W�`��P�jA�I*�,h	���G�^*�W\��;'��3������``)f4�?�or�W�u��%�{=/}��~�6�B��I=�>���hY��t	�^n$����[�#X7��c˥u�c���l��=F��O�Ⱥ�cg�3�86�jJ�O5��H�DZa��hVqʳ��]��VB��c�xe�Fayt"-�����L�5��r9���3G�a);fF����G�ء�ˁ]녃%�u���5N%)�?r����q���Ke;Q�����pr��"1���"�2�"ƃ]�Y]̿���*VCp�N��H�փ���E!+!�+�����hc�I+�~ϯ�e��-�P�Y���O��Z�p �et�Y �9_ׅ8�
CU��D��}݈��蓩�����M�B4v�;/+�]�)�N�-��������-I����>L�0¢����S�x�qgSw�gY�h��^���ɋ�­F�}"�3-�����=c����N�B}'{�K��b�+��ϥ���ق�{�SCe �ˠe7qB&�vj�j�������+D�9��j(�)�[�t�*F U���8 iLh\$k���m���C�V�ܟ��%��/� �9�]���qN����	B/�g5���d$f�����C܋ �!��m9xPE�(	0�����Y�^�E.�a������L�j���|���J��y��Ҡ��Ӓ~�5�
�A�vd��%}�4�R���-��dko�S�7�ʹ�v7&�g̸į."� 88�c;95|&J���@h�09����+)��0*`K]�Tk&�A��ɺZ�ȁ9����l�'���L�c�l5��_���8hw����a�㔽���z�$�n"ޑ����x���������>�~y����_Q���R��lt�y�\��xd�K�G�ʄ�NB��2+�Y���R�$ȟ��eK����9+��l�\OC�������iK��	�Y�]yĭ%	�L���2k���dATn�eW7������N�k���C��}mV�d�ps�P)d�QI+���>�h�C��t5K��D�׻�$�5��1��W(9[ɶ�g5��/]�䀽��	��������!�-�f�Mwx���4��jt��GX��%����v�^�	��_'6��[b�%r�%���U+~%ӥ�
I��b�7��YvY5���of�^����(V3�/~��7��m���({�m�d�����O���3��&�@���jAx!j�lBG�8a���I�ɭz�&,�2.ya����0��������%⭸������L7O\�x�N�3�P�`$4����%}:0Տ�u��i�[oA(���/J	x�t��N�4>�3�u
�R��tc)��c/ҤƸ�oߗ@��_S'��-�a0=�q�y���3��u��-v)��V���vi!$��W"j��ѩ�nu�̏n���@����SB�'�N#�Ze!��*�L�����6�
��?8E_��w��l���R�&������&¤J�N��;�O)�,�i�r��:Qw�/S�ii87��qV�!I���@�o�&�$+�w�}��5���^U:�L��������+[���o�sܗr��B��u�4�u�Zg�԰���!����S�>�w�!��I�Ǿ����Mjv�rg�Jd��K�,VxӺ#��.������O֪0l! ��*d�����8g�3�;J�ܵ,W���F6��;�lTM�d��J%��H�� �f��%Ax�$y	�=��fQ�J�{˱XKV���Q�?�Ú~ouW;*A��Z`Aq�7�@Ay�e2��Lq덊�goB���3="��g:
���4�{�Ե��{�ŧ�i�Q��d����=a�p'4 ��PA��u�_W�G�� �ǟٶ���h絯nH��8,(q�x�cv���=
�)-�o��!4��M۲��u�m���s��)4B�N�>�V������c�[W��a\��4pr��G��`� ��2W�Bj�Gl�K��w�鴨:J�5eO� 0Q�v\�"�?hwXꀠ��Dl�=�ew����BL9�����Y.g��C�1z�C���0��$L�S��T�F��4^8Y�ZQڿ˿���b�X�#��fG�lR���׼yY��C&�@�!:�V�����Y�Q��5p�N)[�>���'�����ca�T�bܧk��Q�����黹Д��^�Rf�Ws�	��O��������c�>8e�~������N:� ��)��7�G^'��E�`n1	�����髲�(l���/2[���sP��jP7�f�L֎��U_��V,�V��h�u�*x����Vw����xA�|H�)U�\2�Y�j�Z@>ۜ��P]_�Q��ga?\|{}F
�Ѧ�����{����5,�s�V�̮O����l���%�jjnZb+]'����nHKI�E�����O��il^c������	�ɇMFO-��r۲�+�Fg��p�6�1p�]��R�sS�TL������p�nJ�/;7=j�,��Ā;C�ea���/����al|�oW��GMH�4<�I7lΤ%y�i�8�K.�c�#Y`�fS��ee=�m&��`)����/������V����F����@��U�1\8F�!6�V|#��i�V��ܙ�
�ko�|P�Q?�x�"�p�50֙��,�S���w��n�Fҳ�ưo�*�O���;JZ���L�6��L*��{vz:qE���FF�a�d��D����H�2���ǌ�Jܯ����`WAm���?^�?��~iY
	SD<]zMg�-{��w��tӴ�)|_��=U��4�u=�cdK������-��[l��V}i�q��T)�I�����xP,t��:>^�c.���vwG3��KdXzc�5�E.O�<#��돕�8k�D�`����1>P��Vt�f|� �����W:�h���ԅ9-�C�)&jB��k�dCT�F�%��!rP���BF�����b6�ߡ�" �3�;U�H��S�� 쎙�w��ۼ����L
���g�̐����V����o���I���:�[?�̿�ܔ+�O�qM~A�^"v�&�U��7wv���I>��ɳwhA��[�H���vG���2s}<�ZFќ�|���,�L;:�W-��W�Q��q^�a��Dg��$��������}�'S,���q2��.q��z��Xq�&���g.�\I�
쌂��u!��R肻`��^�$�n�˔�!ʞ!���3E`���"�x���9|��?�l��d�пX�O[�<��ֈǼ�靀g�2Ln
�U�Ϋ�~N�@�'�u����D���Q���q���;ȭ�Ī����5��ۊ#�Il~=�/(MntK&h�K"dT,���U�2#����G��w�jG�V�_Qe�74&��7�(N=�����*P������
�#�:��
A�Z]G���C5͍:.7�YY��P.$H^/�3& �_!�\�w��˱}O���}��p?�"��;:�?�캷l�=i���))�d['r����#�����m������pї�s�4��]g��*68�k��W��a�DN�L�Wq���Y�9��됤�3�f{DƔo�`�GVja=r�㺔���� ���0��/P®�v���x�"���|7����Os�f?��!b�h9B�ӓ��y�jK��XIrm)8֧���Ǌ����K�x�Se)�J���n�P�P� �)���k ������+�G8���/<�2�x�S��8@��ue-�+θv�l�Ϫ��1��?_�BQSȅᷝ ]�g��[��o�(s�@P��ȑ���, x��G�����Ŋ�9�պ��\|���� 1�('�{X삄���1IO1,r{���KW����0�̕�_�[������hd�I�fa ˧��5�5y�D�k�!���'��C��:��9��@�G�S<c�����;��������H��Hb�E0z	c�9����KV�:�R[fl�qw���:��_�i�n��������7����	Թ���8NX0'���Q�J�5 �$+�w�U�=�K��a�8p:�����W�U�9#����f��SW��QJ����^�G��ɽ!J�_v��:7t3=���=�N��n�〲�tyL��r�/ ��u-'�zV*�{�t��k?�,F*����9�Z�� �9_]�%�2_X� #�z~�%ȏ�b��,b�>�� Y����G�92�!�?	��J�>dY����ڊ�]�Ju�"��vd��z�]_�ۀhl��w}&7P?�W}��_��8g��
i��FIY\��Xrp�[ ��eW��d�0��Xv[�J^C�8Y71�"6P�F
��^"s=�1-��\�Ksھ_d�����뭢̴�K~l�mu{N�9#=���ʴa����u��y.~k��-Rq�7�*o�� B{G��nW���pZQ�����K�1~�f���ww�B��_����婚��W����Q��S���"�n0X���Ьm�}1�gM�FC�
Brq�|���*���D%Q�I��s����G��`�� ������jPDD�t}���q}K�����x���Z{g@sU�����Q������Gzb뒰�f�	�@{�:�k�J]��)�1�zx�Ρ0"w�u�{�!��sԏ_2��v>Hw������}}!Z����o2�����-~��kb��м�D�9��y �����BG��?�����)���gb�/�nc�U:}�h��Kފ]�}�U�s4�0>^މ��W&���G}��r��S.jf���Jh=b�����'�Ha�e�"o�����N<Z*.j��n�3�A������X��[����$�;1��]ɜt��Y���R3.Zm1>�؜�4����*�.�������~C��Bڪn�W2W���s�2���1jA#�"��:<��Ώ�y�oh�~�L?ֳ�PP����k�ՠ�6-�9(�G%.�hj�dL�H�T�GMVTf�Ք=B9ཤ|�QדN��L�����vY'Dܭ����T� �|E��DAh8N���g��P�Z�9RL)��D��/�m��������'�ƣ]� j���U��C�+���
��
L��TI��BZ�G%	�c�%�r}4�Ǧ�݅�����߾=	�Lt��S�ƭ矘��[�+���q'ExM|	�]�Y�b�c�ȓ`0M���KhA\ء�Q�=7b��$7�u"D$�)=#�c��X��f Kt��<�!r�Z�LsLna���>ڪ;���9H�?�d˝���3cx7�q͒ڄަv��o�tB�)���+�� ��JI��R�fg-y>�+��S�L�7��i5���"8C��7�8m�?K����^ᗆ��}��p�"p{���Z/Uͬ���L$����f�?���eu��HQ͋_Ő `z�k�?\���h�:��[G�Sp���m�/���܊�S��'^M}�$#��D����ӾȖ��8���U�x81�J��ه��%9��R�^���~p�'m�?�v������7��z����*& �9d��xEd)oC���@t`:��GgR؏d����X��Y�l��J1/K����y�%&z0���;!���Æq�Ǉ���z�+0X@��ϱ�����Ǡ4	@@�����H�ouQH��>}:Z!YO��¡���٭���}�@ʉ�7_�&k�	�Rާ�����=��Jns�e/3'���Yho�GN�^T�g�$�h��ijY��-�SO��U�B-��3����N�A�F�c�H�,�ֿ�"���o:�a+�o�%��֍��N�n@����]�4��~ş�B����%EY�?�T��x
�]�8~��w��Y���kgO�%&S:�=�@��R�Ç�e>�s�%�S�rcݣ%-<�H�0V��?���0�8ӣ�-۰��g����Gr��i4�����w�W�<#c�>��#f^Y�[8l�W�(`��g�2�9��_���} �N��`�{yb1p�^�Z�C��'����tN���ی.��������b���c��!H�US���'��F0Ɇ�'�������&��$������s�sR�o�ϐ��W�67c���<&�zH�@�фl>#Hwܖ��El;���� ��-�$�H]|~W��$��<�.(��f]OKߛ.;�f�� ϲ3��r�A��o%����2�˞�àE��\K���Ч�+f��ğ��D�qQ��#���4������(��M�'�u�a�^��#i��gMM�����y�(Ȟ#��^����ȼ��#;ZٔV��(�g/���׏G��(��uz�r�v�2<j��BӸ;�h ��[�V��(dC��C0ܔ6@޽'3pF���s%������	8K|�b��6�O��#��B���sy����/��懎c��h���g�g�{~��|+ϥU�/3U`y�.<Q�>I6���z�.��@����cTb��cD ��^Ԋ�_��{�ښ�g���HR��V%�g�u��7���L�;���I�bD��'����ժu[�g�࡜m�ެ�c��U|�e6��s��ng�u�:ׁ�G5�v�=�I�4%/~��dkXvit����P/�`��f�\�d.���h���ϑ�W��!	L���	��5T� �����{�펕n�y�Q�(�T��M��Qc!���=Uts((MQ���������.��4�$7�I���>m��1!�6�U�_�Lb&*j��F�{�X�<�D}�.WW1V�H�����]�Q�=�2lw�6��DJ��J��C���}S~�K'm!��dd��\�S������[w�5���!�҅�~��\����psL�Ʌ�^���d�$��d��B�?�yI�a��d&��6�����r4,S����,�:�,�����M�9���x_��^���5æ�ޞ_#�)<g���PU���.˒n{="gV�Q.���/��JS#�D�r�N���ѥ�����:�l��4��[�~���t2Zn��KVD̠]��b�,����kş���0�Rz�j���/(94�(Ԏ��(�� w_22�3(��>�φ���FSJ�H<�TC�E�R�E?)�Qj���)����}q����ҳ�_��M{	�S�x(�(���B(,����?^�(���i9���<���=�^�l�6�h����܀�X}M2n=.<����뺫���I�U���~S~��M��R|��d�M;�9�H!b�~���g�şȾ�*[��
ԙ��@���:����t�o%���q7����~$Bn-�!�wh���^�vФQ�	g*%��IS;y���<N�KE�!�[	1@'$*�n���g��펑u��抂3yX����mv�K�:�U1�Q�k	�3Kn�f�L�Vy�Hv`�T�,��gEʸ#��~�-`z4�7�*8QhJ�1�zk��WS0���{L���-�Î>Ő>v=ॅ�8���BAy���2NBݺϺ?~^�S��޼���4��5���V+7�ܞ�-U���|���^ʣ��"d����`��0*�?���˾ֵ��	-�(��0�� d��R��?4I�@��J, O,i�:,�#�Dn�"L~o\� G�^���;�֤3Q�y|�Ŕ��e̴���H�\Y&7��^I���|o@����vq�3TJ�]�O`>IX��y�T��D8�%��V��i���A���sÐ�Uw��WTg�m=�s�c�˥�BDu	���';q�*�&��J��x*�C�@�� �VË��op�Xy)���Ja�E����<O\+���ݢ����؍̎�*|*r,r��w��.���Zs��q�h����QxZ�P�aT��h�f���N�'Ǟ4�Y	!�� ^}����6� �cd�X����q��P��l0��� H�頒2q�Op�Î�H"��6PfǠ��r6�w�� �Fb�x�!ݛYo�q(�m�Ai7�b/	�j��E�ZI��h�����3E��}�릊�uXm$-%�`k��N���XI���"��$�.IjYxk2�G�>i���nv�\��������?� �F[�C`=`�i�M~}�ו����P��H�����T0�#��Ǳ�� (����hu�'�'��D8�
��6)Fq��Ȁ�9��ũ�,���2��k�Z*���gl�9f�4��(�S���£;9>�k{��x��n��m�]�=>�����].�ym�|7��t)Jx&��2�L�'�"���+�c�D�U�S���i/�G���[g�.�1� t&��qg�t1zcN12�r�g��T֥�(��3Q���_�Q���^X�D?v�%�-2�j�9a|xڤp��4R��2�ѽC0G�f0ވ��
%|dw��j��ɔA
�z�/Q�J�J��8�:+�P��ǂ�&�;7��
���U@�Z�6��g⏚G� SߴG|��'���l6Y��)��,V��b<@`)�|��jeS�uT����l{�M����Ӧ�g��S������4�5a~��=n���
�'�/驭/j�,ɲ��
���`ޝ�`6�[ҧ=�An���Гc#F�zB�4��g�N���)�ReRKߥ��$��u���ʁn� �0�Tl�곘k�o6V�SzQ��M��+�:�᠔$t�Q�k��u��X��^��nq-]/���� 4X����d[y"ɜn�K� ��������~�
��RD�%�"��6�Z>[�9;��x��m��y����G��[���r�1�"N�^�{��E�R��U��L�Y��N)Ј�s�-5iޛ:�}5F!U�$j#��f�Do
��=W��)�q�d�����tK�v��`���[Y�\�� z�$P>a\�Yo�cN� aw�@�Ѓ�D�9,�Kӹ;p
>��ɿ����ȑ�}Nԏ��A��<���n��jh�u�Z�.\k�Y$98,�z�\E�iekN0<x���sf� \�m %��TZH{��d�`�!��k�+H��6�Sa��kC:��L�P�;Z(T� W��ȓ �����sv�H�=QM0�[��ӯZ�-�[a���!sA1�.m�#IL�;�&�;q�E�b(�f����t6Ŋ����Im�/��D�-�N�:�}��bT��Y�a^�$؏���C����e�P�LE�&B�Hk���[�D���_���0��9jh�te<��¾ .1F�&����J����]��\G�ؿ!4vTk��{�4��*�{�~�/b�	�D�,�g���̇��"�q�"����llz.��sp�%^�̸#0zL-K������^��y���"u�6��N���d6(�ؘ��>&`|0�(h��l�ӑ$t~o�*�P){4AZ69܂�|��C��X56�
�L��l
���IM�vJ�'�8�ڛ�1�t�v���@�X�5X05��嬥Rp)�f�^���)�ZS���!\1m���P�1<f��&��*��lH.�a0pZD�)�şe�/�=�gL�utMo��/*4(�d d��jFQ��.{��޿}y��H��zZq�9�`�w��S��wlii���7�4q�J��0�e�Øc�����ۓ"U��6��F�[i�1���j���m�F#��$Yܱ�,q\X�o]��!�`8:�|����y���y�y��������'#WCU�<��=n몞'Y�4�Q?N�Z���V�����ɱ�J�7;��z��\o�
3������Ͽ|���Y�
졓�YY���\��K��7J�r'KW���/�}�u��E��{6��p[?.ry��r�%Z���� ͭ\d;����yZ��C> �Xo�|�ɥ��c�0��~���
ÌI2r�MBH4�,�\^k��)�ņ��IʥdD.(v_:Pt��2
wj@w_B`j�A6��14t+�˾���c�`�]�/Bފ��o(w�G.�tW�b���Ჸΐ!m!�E�a��/mb�]�G�qr�t$.Ǡ�_�h��ά(9�U�ep
T�G��Y�A��|*�]�6O�u���gӈ�=���X�Ɉ.=`� ��Oks{B���1��V�ջ��;�kV���_Λ�W�� 5jn*)�'c©M,�՜����o+,�&�K��|]G�'�?>�\��Gf�gb
#�v�9�����Εq���q�HG%R�z��]*Κ�Ӵ�!�2Y���k�78�%J\��F:�R�;{:��o�b8����X�K__4��f���ef};��'c�о8ӉS�8؏�DP�^�AI ׆�Ӗ|%�1��X���x�+�-/'w�MUaSƸz¥��>ڴH���Lh$��k
Ŕa]{9��j�3?�i,c����2���t��α1�y��Ǒ)MJh��ƭ�pS����Z;9J��@����������}�?�'P��PV��S�]�чR��Ćt���s�����K��!��;%��K������gU�ϧ���X��9�Mvv�x�͝�0]����&��P2�J��Ԓ��Ǚ���	�0�,��sQOx �����f$-�o��*��O��9�h\k����t��ި&di�eg����/C}�(�R��z��U|�O�(8 �w��Ac��+�\ߞ+O��ܓ��ѧ��e� ����/��G!=%>R��$���Wrh[�	����1>��bIP)/a�͡�Tԟ��CI�(�d�g����ԗ��b!�2wĿ4t|��FNc阐�����Ul�?����|�kHx	Rr��kA���g_N�^ʊ1(S�{W?�Maw�9��|�P�W��4?`�*��I�u�@>0]H�O�DdZ�i�h�_6����O5���(���d'�Vt�B��l�<��S��d��X��)�`��6��I5�'��~���k�F��U�fQ��R�p���;b37�Ts(Bޚ��Id|��B� `V��cB�цn1���Uz1��d�������X�o��y�U�|�F*�O#� O6��~�Q6�0Z~?�8��8��v�ɍ�-�]a��3P��RX�����Ok-'J�I&�g��^OpCgM{E'��*	�ֽ�"PS���(�Y�O��	C����ޝ��U�d�$�a�!'�l?�n��`�4�dkE�>A�p����0?q�M�$���Ro�q����ob~W~�s��R7�Ve�C=J�l��a^��V`I̯׋�'	��72���b��l5��o޻���܇o�u�u���q'�Ug��Cv�uǵ�@6�ٹnR�-O�$��Rk�\kW3̵{`P;U�Bwp�X,��bB�.���Wz�QV�A��_m=W������p:�-��M4�رj��z2M֤^�z�ڼq���¤ه'��x6g�E�Y�l0��~�;mR�C�~;���C��O�W#ڻ�{���|�����i�H� ^q��ߘDתk�~�>�U��5�g�G��J}z@�e�_7�j���j�F�������8oY'q/����>:(�~��	��ݢ� ��;�Pw��e���hTi!W`g��v�;�Dg7�^a����Qe˺�f.�����GL D
q�F���L��h��h��_�gv������;�>��c� ����U�3n樂y�D3%�\��.�pM[�Jm=�?M%	��t��i�2�zުswx�o���a� �;m��BOC�*�6��h���*k(�	���3|�����/���\n�t�r1�(,���W	K��K=g`xq������e1y���wH�������a1G�LhX�ݓ��1�ke� ��і��N����c!���R����C�c�#9F��H�
2�/2H��[K�#�ol���]�6*0��42�b�SCgV� I�����1���RX/�	uY��֊�#d�!�X+�>��f�1��>#��k0����x<v�nQ��-�댕Z�����.5��3#�h��8��U��eu�M��w��'�_�gj>��!����t�^&���S����Ҝ�ց�Ʊ�a5�5)lVXbCԱȏ&P�ӹw=�^?��?�Cg��3�j�v�Ӓ�E�)(��g�|\�N�5<�މ=^����K�Y��yYmWa֓o0���
X�m�L�v�z����ݬ~�O�f�xTs*�g�c#���]Z敳�^��:���j�%�������록`�<HBR��QB���	����VJ����J�x`o���{��X9j>/?C�����k���egє���,�t�O�m�g���U*/j�"m�)�Z��g�����@�B���:�(�u��F���\�m��?�o�u�F��݌� 
d[�E���f���uB�i�!�[�
|>p��<�=	�b<eb�~B��R�r���H�����P����|�y>�V=o��U��5�6�<U
�$@���rrʢ#\f��%�})�;X�����N]L��n���ÉI�fd��+�v�d���&�Vq�
'��j-m��q+"��wFߓC�v~b�v�Ta�5��*�'��>_�?�o�.W���I�<�n�����,`fN!��=X��� _.31��#ᘊ�?�O��A���.��mF?�������k�� |>�>���c�$�����(��A����励ƃ����J����⾗CUiE�j!\�����?��!g:�-2��XR�>}27�����Z�+���D!���%��m4'c5���~HUO�ň-�D�ƁC�(�/'�d��O'�RIx%��-�"f��!1֫z�\]eo�`�j��k`�IXf" W�U�C�n���w\|+����GB^R�t8�麮���dP�~�����a�����.5�������➕T �z�]��C��t��jT[�dj��R���� 1zx���V�;�Wn͇&�x2��R��I�E&yjp`����=�8��B���L������}``9�4��#Np0w��eg&�R�m�or&Q/�ަ��U	O�!�>�	!%c86���[�@�f�~T�r�Ā^:��� F�o����I�l��xoI���R��(��DbD����x��;��ު9���s����W0g@�c���jZ���E1**�*R�a����l��<�ʂ�7Ƥ1}�އ%S�(X���d�+1�_�5ə䠴��Nd�PPX�)M]���>�4�[۟�&�M�(ݝ��M�+���K����[Y���}������ˆI��?��K˞�@gu�ߨ����nŔ�&�=QU�3�#�{a̹�n���C�_�$J�ǁ��m73izI�yaݕ���h�l�|���	x2Ąk��qol���)�j	l�og��u
��C �z���V��WO�^|&'���c+p�;H˱�ȅ�t@5��+!'���@�;?(O��4�dl1j��2�m��J!� �
F��w�("�K�
pƖ�LK��R9�S1X[��g�s��-&�G�KV��G�3D2o����zHa6�Uj:z	k4���j��)�!-H�rDX�B���_6Zp�FA?~,�,�z����ݐ�t)5Y��!Zg���_z�f�(���{�?c9a�W�̻���h ��
灞��v � �ˡ?���F�W��zz)��v�?%F��RiQLU���)6��|�t�j�!�t��yy��E��m���?��(�41��n(|�3�tUם귃���䪰�4�+\U��������l��[�1"�<UGi���f�����>>��*!Qm�<+e�@�����qsY��T�����t=q���y�@�)�%묓jw�.O�(�c���.�s~tT��<��	+se�('fi�^q�g%ǟ��ؓy/�	���~�ٓϬIo:"B��~�C ܂�d7�}����W��~���6|�̗��߫G�O��/�:3�!+�~Py�	�4.�y�n~��h�ǝN�Gɚ�p��c��21�0���g�u�垽uqu�h?/F���.LC��~�uqzǍD\{�
�_�\MD�s�qO>�׈녟B��Jk
���/���w���T�Ó�}�������e��y��U1��g�k8Zf��"�o}����c��Zj�T��R}�ٍj��8%f��/N����\�IX�i��ۘ��Z��73朆/-�,�^�kcW%��sS?�u���9�1�ƚ{i�0��\�[Ӌ��hᇪ����z��	1N���$ޛ�Ev]����3�tE pZ���|��X�7΁{��f�C��Ό�/�ǔ�ߨ+��������@�QD1����k\eaG��k����6Ke�k�c����
�� ���A�f��ǥ:6��W>�|y;������1�gkzq�Z�3�qC�h�]�v�_�.
�²��[d�W�w�r�Z�������e3H(X�+��K�:ȧ�P�I�(�