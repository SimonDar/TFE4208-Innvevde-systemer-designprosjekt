��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U@W~z,r#���7��:Ǻ��Ƚ9Rپ�����91*F����Aj�!w�Z�O@��A�u�a�$�"+Ta�kX,F��+�R�M�-�d��T镹 ��
do�V�b��
s�9H������hˋC+>&�a	�� W��+n��;9:rs�ա�uۨ�N����n�x��$�z�]����)��7���\��ě*���y����F,f�=�4p�}H�Y��f��fM���u�����{_�w��۴�;�iKZp%�|7E50�`�wr���}�����'���V݉=2�5��Դ�^��ɟ�'��31݀Cj�zyH#�{X��놳��c�|b�[��>�d/�YQR��k��:z �.C�.q#W���_�F����O�Yf<U�v	���R��!hh��c�B�����Y>�ō"�zBP�w3�	�{�*�\͸��V�F��L���9d�����-�`��t�żV���0���2��X�XcV��QctFF�=&	O{����#/�)���H�S����1	��v�7�{�<Քh��-����>%�k�`��`�Su����|ׯ��Z�'�bb�)�ܕ����o[m�i ���{�4�3�^�~A��yCL���_��y��H�{d����O2�������1TP3�	H��ʣ�{�k�N�j���;ݢv5����4W��H�������DH��5��Ґ�|�~��~ܭ#Խ�A���.7v[�n���Ɠ6����ʲ�J�2;'a�t��E�, p�I����y�}?�b�U�^d������b e�\;N�^bHg3R�u"��������QI3�{�n��.��2��ud���)*г���)�Dgb$n|�N�jҁ����(���q�ɾ�'0�/�ᚐ_,������hY��{������W�х� J.|�sE�"�!��$o޴�gӡ�SW�>㵛E ����ZT԰������<�L�-`PV��x�C��������Є���9�����>����������{�%S��t�T;���!#�KʔwD�fV�c�N_$�R�F���hG�?�[�"�����4��V<W�ԼgЁ�)���> �YF���z���t��_m����QM� ���(\�)�w@U����.�O�K�;OKs�G[Bx�����@g{���sL1��}<6�n�~$54���U���s��m���l֫��:�ZG�{1y�u:��Q0y"ָ:�5��d���9~1fI�Y�}����Eذ(����h���B����h�a㑜'�??������r�Q��,�VJ�����V��������{�� �hT�H*�7�X8_����-�R�׫����^�M��RM��υY+r��	�/�k?g����'灦
G�U���L�$\��/rf�\u��2k��z4$"O�~��|F�r�!���Y�n��#�ǖmцQ��Rw���n��?%�(_�ځ���.��$�_�1����|ȿ)��P���S���,D�+ri̸{ֆsT���u�[�Pmӈ���o��%S"GZ�a�����&:�
���x�ZD�� ,�6:�A#� F-�+K��O���a6��jV�-�����ޏ&\{ށ	P����	�n(��po�P�n����[@���E��7)�'[���t���B�������j��7/KB�5N �fR�1�v$JJ� �筬�̈́�<��4�J����{ ��{(F����_Y�~�oa�a��+��F�j��cc��~�����4@-Mr"r���QȾu�;�pA�Pg#�~n���(��b|�~U%����������%�n��ÍfzՀ�4s�F�l����ߧ� ���P���D�Օ8�;�7�OJ ���*�!No���8!)xX◹H($f��Y��t_��P�J�/�Z��ㆪ�ۧY�qd�r����F��o����5�& $�wUڗ�A�St�M��A;3���"�Fxʴ�<�Gw��,��9���p�m�p��B� ic����S��(�X�
D^уO���}�-q��,s�l��"wϤ����Wk����?�A��72H��WF���ۂR�����m�z�����`(�g^�-=}��{q?qR��:���y;�)u����95(��eS� ��TeU��_M[��WQ�4�A:����Q�NA�U؄	�[�P7�q��v9\��J�4�l'h#х�Z�s{��/1�GՄ]�J�C���<� p���g�L��*l*�L�;s�C7&R�픅'Qv��2
����F�ȩQ0���,g���\�W/;�'�=�PmD����gU��b^�j�>��>� �L�:rݱ� �!Q���'�03PR�狽`�����ޘ�к��Tv,n�\�=�5���z#�O�BT������[[�~6�*��1��x
�Y�q�^�zxQI�����r9�uf�H��	`��PH�\�,ͯ���[p+�n�N�~�����?,KW-���/�%�*!?�)��r��M��A=���l�����#��Xzt��2o�L��ZiO�ɶ���ի�wG6����Q�N�����u
�&1��#�I	 �0��z�$���_v���\+MWo�5�7`G/F�S�s݅�g&�x0�j��.Xߎ���\Å� 2X�rnQ�aI���Dݝ���_���|�c�u>Q��n{��Cw�������Ⱦڅ�'d��8ܭ\����7׎)�lϝ?q6����y���	\��2�KCf���׶�����9��0XlM�^n�d���B�h�v����7.4�y>�g!�#�a-ѾIV
��8vOf�.��4?Ň���5ێjor-az�_��6O�ZeeƇ췶�SZ�����J(���x�]�YV�1.%��B^O�O�����K��-�09g�/�M�����%�䝺�������A�G�$%)Y�`Ҵ�M���@��(	�a��v�z!����ݸ^`pl?$<�{wg	�7!���:�\�w5��A:~K�<a���[E2�\j�|��IU��5LLr7�>����I���նy ����Y�3��Sy��O4�2�y�,}1p7��L���m��e�(��ώ2��xoq�v:0Ǘ&�A��}h��˼�d���q/��#͍���/���X�w�8�G�F,�ۿRӕ��.ʮӜ�9��z{���z���}��ɖ�(�Z�X1���|��o:-�p��
ˡi��D'��"!��D������r�ŢR��g7ľ���*z�Qi
�΃xϘV��x"�����h���<���Wi��@�`HA��v@���v�����V��
"Ù ��/�љ.�ӂT�ֿo/P�/
�Aq@
��Jp��5�o�T�|��l�Mě��Y�E��p�`��l��4�I0�ZB^�`�3�w2�s����MjӪ���"�'�0o�Mp'�k�"7��c���sO#�X0��H��]�Dr3�<�r	��Q4a�\��ךSY�v%�Ƌ���SJ(�1�2+*�!����ϐ��8$��@��Y��ǹh�^5���-~���򎝾�l\�;G	mVvφ��WQ	���j�	���,z����n+�X#E>�R�TA;�Ӯ���,-�Z8�;��ɋG���1���x��aHyh��ϓ2��+d����)^�WT��=�=��}�M�2��b*C:Ȯ�/��|���,Ǎ�Ul��W�[�1���Q�	�/*����f�����j۰�"�C���?�O��n��8NHr���"[��A�*5�ٛ��oͧ��^g�e���%5!JX+L�c`*w�Iy{k��`���$k�W.R�Vv�sُy����I�l���%�*\��ڥ p�5&��8I�`�x��`�ldx�Bb�p̓p�6�+������Z��G��*B _q��p^۸��㳐hUڔ�⊉,�Ů=3�*l��^�[X�=K
�b��)F�j�V	-�ʝt�y~xi 	;�t��nR:��~FbW�Af~�
�!aq��l���7Z�ƣH�7�%��I��wS.��[v$�ŵ\y����P�
��b���H6���W6�GR��̈�K�I�eYة� �E�1lx-':���[���R5���%�s��>b
�H�;��x쾎1HIGhcz�� 8J6'�հ�?�Z�u��N7�'ܳl�& Z����=Xf�s@w�V��YȬS�-��
^o�#���)�^�O��P��`]��8���Ὼ 	�0/�Խ<x��� .^Q�%�h�|<�������+��2�6!�����yb��U˹5m��dл;QL��Ƹ�\3$'d_�;�� ���0����8]_v�wd�x��4��=�(v�-+CN@V�@\�ϵV����z#I�)�E�%s+ �ڎ30_��%���%�S����W�����gڵ�l�)^Q����]=q�h]Z�4,'"v3��Kz��1�H�X�\sl>��v��R�×��6��E��5<xk�+MA����*��kzU ��8�񤙄͛/�4� r��%�csw��'�J��R$��g�4���[Ϟ_׉�YBn8����X!4e�b�M�(O�V�9���rgVQ� F��,�P��Oa��3��R��D���ݍZA���\)�H���(\�����t�I8^p3Xs�c���mD���"���pnl���,9�����H%�D��G����hoKAs���po�p#ˈ�5��QL?R諜q$��P7�b�7Yʼ��Q�8n;V�v��+�{G�"=��@�Y�Õ3Y'#�V�����b 1���-N<�ɓ9�&�D�~��v�Zj@X:X�0f�О���#Bhϊ|��Y|#ʮT��M!x)�-u��/-+]�=����3j	aVK��tk}:5)�H�b�NQ�6���4{��Ő���
���M�Uf9XhUk[���j�~_�ڭ��b C��i�3]�f7]0�������IT��녖���8HoKr.�����K�}Y+��É=���d7���Y�U�񮄓8�Xr�}�zu	��회.R�X|I�gm9�==��b����V�׶|a�M�?��:���|l
�<
�;�n�J���5w�>�|,{��Mы<�)q�ia�m>��K�9�Ml�bޞ+s0]"!l#`IC�D��ѫ6?� ��Ld!��*�Z�9l?�j�:\�ЦO7���so�Ax��n��f���ފ��OU�ʘ�>��Ϲ]�J$Ss�/�/霑�NS��9Pt���fh��[� �U5��jB}��*�Pl��t�,��M�K������Fuؤ���E�r{K��d����)10Ðةo����I�l�s�Ih����:E�@_j��-�K�ES��5�}� m$I�V�s;	�:�p>�=5��El�#bOC=���O-y��
e��&=��|s�@p���U����3���O��,庫Y�q���M�[N��`7(�̔�;�面�L�ʡ�洞P
�;����ΊZ�m�Qj�G�Ԁ����~��V5�Ӣ?����5mR��j�و�ho�"�Seܕ%˹ ���;N@��l��^�������TU���T4O%_N~�Q�-��6�猏gHm6�[�G�c��.S��5�C��/V�O>^g��p��s���d��$�_��~@���C��� �
��yT5#9�_{�Z5�	��O:G��n�}�p
�Ǿ��.�㩉p~Ôs7P��a�M�������p��rףe�b�2�P��HȞ�r���]�S�{#��g�Y��/� ��pM�Zðp��@���K	epHC���s��;N �@�b�ok*�G*�dP�����Ǎ�SR^����6�pI����%I�}ǋ8\EHrV�J�����Cu�xQ����_�(�)E1���j��[B�������mY����s�1h1�?^��j���s�m� �����C�'���P^��l��*�H�u�.�h�.SdK�~<h���+�)=���[qA�/TE��M��ҝ�'�"�cE���rFb���p�Ae�@p��H�h{%ҫ:��؛�=e�[�Zgŧ漦�A�I��s���z3n�v���6J�a�]�з1��0�M˲�+�q7��Wn���!��s����\�9T���P�$,X��YhkJ"ɸ�v�j�����E��[p���� �*��sJ���D/7�[�kYow"6�q�6�]o<�&�9x^�5,r�~i%�H��wX�|����8��! L���|�l��vݥ���i]f��^WFP�t�tj?|774��W_���Ui��wZR��D��8C��=!�l���o̕�B�K����˺�z�D�k��%�>�,�I*�ɬs%��$)��$�xR9��:�
.'���G<�ӔpPi�a��~�P�s�����;�ϳ����.M�PU�c�QKo!m��-�p���[�:�S��9Ef�O �?��H�v�.L�E9Q_���8�J�d��ė��x��M�"����Q-�x[7k}�c�����p�}��s/-fĚi;J���r#@JÊ��o��/}]Z~�.���+�AǑ�l�u�5ny!O�*�����s�[�=~��aT�O��0�(��?�K��{�R
Ck�������%7/b��l�*%c�`�R�O�g���f���Y���Q�3�qȔB��4�H��f�x�~�j��V��������(��n����1P?GW���e�w�%K�(��9!]ƵB�s��H��F��"HEx�{䚈oܕ�Q����#O>ȭ+��eykj��j!?���j�8��:?��Cp �Elz�s�a����]���N���r;����&�^��[ƀ��
���2BOuX��hW�˼%M������8)�g�è��)�y��J��1���\�Uz�h�yՑ�4{���F[���xY����GX��ĳ�E0�S���ǎii��X�.�g���7snߛ�F'���y`�j�����Pa��L;)*�I*�;�km'�@XӋPu�ahB#���;��p�\�
:m�}a���I���a(�n3�����ݩ��P|Þ�Z��Y�OZ��1f	%I�K�v�U����q��w���~UX���gV+���S�[(\��KY���`��L�R#׀�'m�	��<
�`�J��&a�(F�%���v+���TC�aC��]AG:�C}Έ��|��6� !��h�����\�Bf,�|�x�72:�+���ӌ���
�*T�s�UO��h�u�ƀj� I{�&�X�Bi���.��0�^ 7���US�ַ���О�$�&b�M?��9Q�ߦv�'����9�^{��I��H����.�]�)��k�<�����s����H�����xN�m�r��k�h��z��8�j�G�|���̀��m�����Һ�0Ӹ�|�4$�pޫ��A�^册�;-�r<��$@�W�3�<G25�\�[�8re��|��QM��iU�-�34��ݼ�ļ���2}��������!�Z�b>��W��`�v<p������P�e��KV.��0e�4yt|�~��ZI����h�^��W��gl]<tx6�kN	������8���[��i�pAd�O�e�w���+�w���A��w��������5�|�̶jD1Y8�o}^�Efc�>��8$D&���Y��3��]��#o�q�Ga'�>������3�O�m���!8�B�0��+��7�:�����X.�����a�;����ڤi������Km��g�������rֳ��p_�X�"��h1+C,e����F�L�+�u�w%�뾞zM�b AĜP)�3�V��妎{v\Q���V�^t455B�Jp�BG �7��w0k�U���˵޸;�T�.���1����<��{&�_�<-ц^!���Kk7�J�!�2�OB��i_ԩ>n���-�XL{�� |���p`Z�zM/���f��tvg�ԨL7���ЏElt*�K-H��e��zo����T��
�r��32x�6u�)�0��*�J��#�$��lm�`Z��w��ivi�p���)��<W�=ʭ�*�{;/d��o�P�T���Xp���Od}R�b͈���P�^>��K��k�{���U���_B�՞�*�U����i�m̟3k	J�0�
�cd`�ԴX�AË�L��=z����>�J>�~����i~a's��Z��y��>u��g����*8�n�m��{=w(���-�o��cJ�@\<{��0��J���름��H�~��d	�5�u���n���:R�`ܸ�³�΄nY��^��k��(k~����M��Z�`箹Cc�<�p����5F_���ұ����va=E���r�CR�D 9�qa��̺"�t+����}��S�u#�9�a�V����A�w��U|�9(�w�	WB��*�
��EUy���(JXo<|1���v�(�xɶ�~Ӯ�h��;�ˇ�[�m�a��@�C�MO��'�d�Ҥ��U�,U$���N���=���Қ��M^t������ň�]��+@��2W�w��]$_��vN\�Z�V���kM	S��3O �v�}�'��mƔ���o�E�^�P,�G���E3*�yA<o�D<�SF�.����Pbk���~��M0@��y�'�Z=�u��p,�oorO�i�(55��ʹ���`r$�:I���s�eXC�|fM�ٟ�u�P�mg�v�!�B?���`���8�qc��㬡�� ��\ (?	2%�U�ʘ�0�_}S��Q?M�IEb��x�M�J�fF���v.�{dA� �'l�ţ~taS:\�|W>c�p<��R���-��`�g�FU�j��G���UM�9^){�+�0r^��Q�9kzn'�Si=!�Gj®�����D�쉞�ƛ���>��!��z:ғE�隝)x:�iά[�DF����:ux�� ^m �`����mkA9�y(�Y$� A���A:G�1�4|�@'�� �J�$V���m�Q� ���7�<|B����Y���gGM�!�I����p�wh�5hM�E�(b���c�/�<fO�ck��V#/׮��&9l��O��zx$?�����|ɶ����.&�,����/&#+ gº>Ya�z�r!B�<,cc]���c5,�Rg�?�r 7۸��C����u0;�F�N=�{�A.(EH�l�lCJ��VB�z��������)�����N;���~����
cX�/y���IQ��}�9�{ֵ�N�J9�ãxϣk��"v��2
]jf�q�%LR�����N��3�PՅCV�˅��u��f�ڌn�N�t=�: H��.�zB���	�j�^���Y��ഴ�9�qU󞧀� w�㧐�g�S%m}���:�|��ݡOk&���R׏|@��R��De�@uf�g�� a��/)gu�]����O�E5�[�x��Y���nK�5�
���Z.&	�!K���n����L��f@=�)����׾R3���/��8چbdt�㣓/� ������`����y��������A�N�B�e(a��a�Q�y8y�G �ߓb&��]�h��s	�\��;WV�e,"d{���Gɽl�&x��!�+"<!�~��(��~����G�wPza�F`Kp�Xu�p���(	�ء��X�w)��ͱ�b�;rAS�a۫ SB�l�3;L��
!4
:6�Z8$ � =<yڟQ�q Ĝ�(};�B�"����:���Fs�־���a�<�!0��z�h'�V���!�%Ϸ���b�-�}6G�����j R(�;�yq����x8����� E���'���#//�u��$a�sA��Z�L����汒{�t{F���I��3
0��S$ �%`َn�N�j� �P;!~S�ǮFL�zZ����w�}��cM�fV��;�����P�b6�0���?t�|"���n��'7Q��7��7���[��Ŭ��|���^�F�@����G�����U��7�t7���*w:���ܡ��(ﰹG�@��Sǒ)����z��O�ǩ�I�Ie��5��{��P���[
��q���ΘA�I��sD�a��GN_�M�5��&�1���w�,6�8��A��$]���ef�����!�cy��{؆|a���^K��۽���1n�?��M�o�5}s �z�z�V�Wx�Z�>��v�Ӈ��pDuX�k �R�t����)ْ�G1�F���C�.�o�~��a{���Yt��Ƨ����7�����g�[r�~1���j����WR����Ɛ�����K������Q������< 2x��������$�����2��	(��W�SZ2�MF��NI��ny���M�1
:@�����fQ �d�ˊ�x�1�2��9a�!07�����.��Ugܣܷ`�fv˄�S!�s]u?���]"?����Q�8�U�%�+�LSJ�̬�{� ��*�B{;���bԹ	11)�1��h;f��R��k
|���\7�m_���,��Tݳ�[,fC���,I��7=����q�o���U-d?��JNY+.���|<Ə&�\�MJ},I��h	�f
R���n���vCƀi���3�������DIm�9o��9�X%[�/ؼ U#kJ��j²�)@�<d�\Mj��JV��ú�&q�[Er�E ���u|����sm�dY�#���A��D��"�vjQ�8`�j��/�RT�=��'��mȊ����)�U��M0���qF@�=C)�i����֭�*+gJҎ���Ǉ�#T��Z;��u�hܚ�H��R]��d0�>�P&=�2i��d�g�iw\���,�78�zd�w��X/`J�E��ğ�;#�	�7Ү	;��F.5C��KoI����#���b��*�d������F�y�v��=��J�ǇJ��B�Fv&X$��D)���=��ƑY~ݑyݪ6����k����F(i��f?�|���/���Q+��Ȁ��Nօf��K�ԜF�zO4)E�A�r��(�L��g_��Ēe��Y'Y}R��K�S�7&�ۓY��$�wAjZ�幆Y��@}��4̴��&@*�����9���4���������qھ:d�3(!���#�s�/��S�S�h(��:H."Ծ�TZ��D�\��Hu��GWy��	2�福&�'7�E��o�v�� ZE��cj�w�g�y����V����\�͙�	���C�$d�-�"a��E��T��������n0��cblI�<2XK����N�J\}Z�e�M�-1�����	�f�3� �!ݎ
�ަ+�t7��XH���#Iųf ����z�����Ƙ������SH�E.k���k�)��Ea�8�	�E#��?L)).2�ɢ*N��u������[�*��f&�;��vĪ�yװ0�B�����n+�#\E��H�w5R ��B΢Gד�>���X��IN�g18F�T�����Z�}�lz:��\��z�j�_z�ţ����{i�Gh��M�o+�2�UǞ1����s�1ud7ݛ��Z`��T��A�'�+��翟Ζ{b*�x�w���`��tH���8mO�y�ks�4�J�4�&Ma�X�{E�K���mv��Y��Rݫq�Z+�����rՖx�G4�
��%v���Ӏ�*G�Jy÷����N���W�����o9��&:&����?�TYM��b���/����w�r8ݞOQWW2�����v�C[��/j�PO��Y:������\i�h��/���t~f��'�hʽ.<&\�ݤ�q�����0I%�:��IM�sC����-��Rk�u�Y�V����Ȳ�����J5�$|����ڝ\��A�)̿W���A{�اK`i��u�q4m�7V��>Xj��:�ů��L�S��z����pp���
Z����o�bs�'��Bxܼf#큠Ln�$��W��n��7@����kM��dy������.�!ƜՔ}3�05#k�0T��I煈M��z�G󄂇o]�^5phU=]���G�To��mR�������"�鋸�+�}�`�zR�����,�?��c1,7ZY |/��/�p_��n���T�	�R���� c�b-fW�$�GŅ�h2&��U����嚤I�`;�b��lևƍ:?��3�r^P��TF��8/����]��h���{�.�,[�@����Z�o��A�Y␍�"��""[�Po �����	ɪ�j*��o�� BPO��ET��t�(�6�7�A M���
����4�e�ߴ�&��Fbz��ڪ�69�'��})	����QO����#����Y=�����K7L<�3|�C��O{0'�:�^��y�E&�n�MR�s����q,é�pwU8��M�#M�ou�U\a�Z�K��%����q���#�^�X�)ʇ��B�0ۙ�rCw*�Υ���N`��aE:�Oyk=Ch!pƗ��.�L�HV�=�QMw4��\���#R�
�S�z�ҺR3����ڧ'�l��Rj�5�1�Qm�f���c܍Q;��2��wo����Ve�{�+����M�	� ���`#� BXQ�L�͠�9���Q����x�q�����*��=�lD��NtLi�6�`V+���8�}����*I�'�������j)�m�SIa�%��haz�.2!�}4�C�;�,;vK����n�������Լ�ڝ���Uά�B^;`v���c�a�\����M ܸ��N�)��w9�$��ZB>��
���K�3W������}A
�?��t\��!�B��ԛ�P����TV���΍��9�{j�M{�M�����q�P|����Qd5)��D/{�S�\�������Z��(�G�����B��}�m�{����C^�,㺽G�x<�5�����v�A����)Ҹ�h{VΘJiY��a����5�l���e��3yѕ�]/?�݅ISڧ���^.����px��r!�<��Bl>��T��6n��M�[	 �lj�<
������3�1��!·�I�%����E�������{X*���B�Cv�EZ,F��-�"�&�<�5�c�gT���u�����b_�]�G�jO��a p�8B�0q���+��Z���$�� �����0�8��ML�<���1A��M;�Rf݂����ô�@��l��LB����I�e���z�g�n~z-�li���@�7T��i���aR�Z�Vwl�+)#)�տ޴ZX�XÑ����>ɷ��>�����U���?��j
A�p�5���Үxp�5��^�i� ���0E0܅���w��ʠ����
�)��Es�qP5�Lf��x� �T�7ؿK�
Xy��1��Eabl�W�3�	n�HI���N;��i��
��^*����7\G��Ǥ�G����R7&�wkf�	�)��Ň���ð�H¾u���G'����.\3Q Eɋ0�����}�W�p�Pɽ�[{��.����&���J����]��y���
`o���zt�ka��r �4��͔�J��o��y��1����@5z���d����!#�����y��ب���'����n��1OZ:��>��}�Ɵ�l���%�$�r �|�Qa���l9`�,'k�������+f
�t�b�R�����Q�X��ј���q��ڸ��<���aŃI�r����ϓh0$���5zy:,��/
�仆7v�O�ү+��μ��B`�YodxJB'���ؖHM< z]y**�����A�O���8�����u/O�4����8'��x�?���<�"\�`��($N���ȣ{����L�-1e�����oӳ���v�d�z�����ɣ�˖�E�9c�,��p���Guӵ��ο�MxZs=O/����ȇ�!�P�8�<����T3����F� =es��d��xӼ�r1��b�>2&����Ć?W�NQ� �q(�T��9u#a�f�_���8{�;��f�+����ȝ�ϟ &g���(|)2�*��2uy�vY�ڒ�}հP_�*F�xG�����K^I���{�?3�����@G�:�2�"/����(l��10����4%�6�0����+	-;�m{����,S4�11�#�r���{�j�'�=)�K�����p��88�)XH��,��݋�����ќ�*g�J��8X�h^ї<���t�`g^���&�ߺ����qN�~��')��c�L�X��E�XK��f�$�)f+4x��.꧉� v�ϵ�9���wغr���d��_��
�D�I�93���S�۱h,��(	mU�7Tޟ÷�4b@�x��Ȇ!�X���+�=Xݸ'�����v�JS�w�Y����I6�I,-�@8��[s��T/C�tY���j�8�L߈*в�p�v�$_>��-��dqA��5`=$�'ץ2�z'��e�<�oJ��l�S��A_����l����N@l���UB}���J�ѯs>��޻r.�s�Ϥ�����0����W�鎯�
�)� �N�UCwc2ΦN��Mg.��7mY�s���?����Ib��*xg�ת 2B7n�J��x��&.�x?�'%<\{�gh��t��:�^w~<2���?ء�d����)f@�{Y����.,/�9�4-a�ä��~�u��zr/�n�4�[R�Nݹv��H�Ә�oÓ�3"ڈZ��Np�Q E����m���̊�n��I��9��T �o�vfryz0x��}JW�I�Ur6�u�@��df
�-�%��3��|�YZ�^�l�&��c�=h���J';���i���D�(7X�m[yj��Å^=R��G�k�.�x�|$��Kc��=?�������)���r:b�W}���MIRL`��O�� K�4C.|�Ҙ+��Xn�����'+����a:ޗ�,��������&��F���"N��x�
jOvj˵��8����qw��H�m��5p�+)������,�����us���v"LT1^kr���p$�����EJ;I���oN�ͷ2� ܷ���ִm�Oa�`W�2�B;��)��rĹ�f�a�QL��9�� pVe�Hh�B��N����}U�y�rx^�cn.]z��g2�H/�u="dT�/��":�
��p*�:��y��z>�MQ�Q�֦	|?Z�=Q���?��j�����Uȍ`������n�?�rc.T�(����z�쑍�Y��W
|}ے��~�rћd\�^�$ђ�X˯S�򲩃|���~��iɪ��Ht�9�!�~ ���6�z��OP�LN鍔��R�����3�0���5���r9Q3(+�=��˱zG�G��ǉ����+�U�W�V�t�C�18�v��3��7xq�7�e@�
\G�4P?��'�� ?O �J'��h�,��X�.���?�+�O��f�X�����!��}�)e��x��SU���L/}&�6�F�2���j�/��;���Bd�i�+[��9��n|YF��k��6,�ٓ6�Q\B�71�cn���t%��-l<�|i�*�����!B�<�oET���y\��_�_��c��_� Z���HP�:JV�
�6{�\.�c,uub��h�����u��G�<1p�۽,ޥ(�S���氤��u"S*6Zj_w�}�[�iF�5�4E���o��{��>�.�x#���h'2��W� �mj��d�� O)<�Fi��/iC��q���S��O6���7*��~w� �Z��'��r*�l	���qb��
�nѨF�xW$��A#��e�5&���e1jό�0��\��B9�'�;s�l/�,�(/&���|[d7�v}�:L��ʄ�t��wpf������2nf;ZP���~�8	S��4���LhY$�lGe6�ӎa�=9�YqOqZ�����z[����h*���I?���E�Hs�}�!5�A%9�ܵNZp�0�KX� �7�lۥ(��Ys��O#�Y*��9!��s����}�5�^b� ��CG�&�N��׃�b��*Y%��bp/8�w
g�A\�^�ڲ�,�����u�-"i,2� ��6;�Qd-�c޴7k�I�[��X��T�SX��S
���C�apt����V��ڰ^k[j[�A3�"$wv�W�d��\e���B����&^��t�r�-�3���ke��U#�,�ߨ	���h�2,��7Q�i����~��I���oF��b$�ՍIx�m�H~W�	�]VҀ����*�X�b_�kXh*g�˘�^Bڨl	[u�wv�,�A��kv��> �!���-Y��5zA��K�6�*2i"���汹��i�����V��Y�"�� �k���!���#
�`�/K}rDNn3p.׍@��uh{7 ����/���qԦ8����t2�&��+
M�[1+wF�YA<&��1��Ħ�]����N���QtDFS�p�pq��,5�^���a	�l�a71�66�坹��z[q=��4�NZ5ҟ�2dȴS������s�p�.	W�{&�{��_��n�+�S�S�zу�*�W��xC eѼ��r�ȿ��Ld�lr9d����-O���1��u;�.5_J7F2.Sg��1�9�1=������>�U����4H�G�b����:���;Imzc�j���XX{��)�?4Z����L�o�ʰB��f)����u���J�㫯!.�-���1�k��Dv�!C��>���H��9G��l*W5>��zs)�!P-����t��{���đ˯�r��
x�
�� �q]�L#YW[e��ܬXct�Y���/֊k�V.�_7ch'ɩ�����bzb{��g���w�Ep�{��C�o�/��7ED�D�����LO:�v�g�N��	���b�����O��ׂߑ��L\@=D� ��S`��Խ�r��9�%ݼ�C��x0�Oh�<�]�Iۢ�D Њ@�p+(�g�*���A.�A��F_yO���٘�kn�m��0�uw�vS~!z80 �@H��� p(0�����@GQ�<��
��d��'�������F�Q���Dw��3��z-헐�YIq�{��.;3�dh��Y�.�=UQ_I�K�to����c=��-ԍk��Zk� �o�����钥��9��@��㹡e��	p2��N������n��><����xڌ�����3���!��*����	����_(��)M�{!$�����P�$7i�^�w+��cn8¨]V
D	�	�&�Yb���,($�k@�k�E�T]�祙���b]���x�����d5��Լ�S�!�l$�=g��N(uL��k���5�_���N�ɺ�6����B��`�|�13�+�q������)�2Jj �WϤ&+����?���\�\.�8�u�F3��)+^��ԎV�)]j�hjMϗ�F�߂���d����4/�_�q��5�/IY�U�-j�Q�7�{Y�g�N�������$�k������|�[����a�����hS�o�ɇ�Ck%Q�u�|M���|���J���`�5]��o m���� ���
�ozs�GZ�L��U͐�!�=s��2�Dq�1�{�x/�����f���\9���y��X�bF���o�s��V�4���յz	�iQBߍ��Q��-�7]/"�x2 e�I1��
YMB�:jzW��g�U$x��ܿ.����5o3�(��,T|��'�LP��k����ۓIp<}\x@���T�Dw�������;�̒�භ���B�Is_+������a��n"u��� �EMRv��נRp���jX@#����"���q7��u/ww��_��V3�|5�tm~��~�S�CS��%�Ob?V��bh$y�g���߿��������w�^�#��4Ȅ� ���h+�'+	>+MkaK;Ar2�9��}�����)�en�2�@�wP�����g@���0��Uh*��;f��]vo�0W*t:�m�����D��8t~x�����RrW?���лi� K(�kI۷�6Oo���vf��L��vԣ=�j��ƯR�-�B��#n�2(&nL~_�+#���M�$"Ƒ!�6�Za����&��|�K[�c0����lE����a�����"#��.Qյ����#%o����k�HN�K�_���TE�;��ij'����~�����ާ�t�F�o ��6<EH�^\[#��(l����� M,�P����,�C�%���s�6^��ݪs1<����g	 A���n�9r���Ü�?�'�A
Q� �"zD��9���.�oi�*��Э񱊹���U~T��L�m�W����j��~/�o3��p�y��g`�����5�2��}�n�$|����!�sw�_�)��b=9���ڏ�5��W�v/v-�}�ɒ�Ov�����W�q?���L�T���������L/*m[�i�?p�Ymc�_���&�c�.��x��[�D����.2��b[*�8-�6�lF����b����K��E��}f����g�h�a����+�����~��4�D>u��bo�H��}�9��ɫT�����a��A�b+�B��E5'u�$���_E��wP��Y͒j�&�ۛ�jk(%>E�H@-�mP����qi�����&��$B���桀9�U/I2zsր���r+㉖��;P�bt�><,��i�h8�J�fZ�&@���v3�g`�Ƃ�^��l�� Cu7�(R��l�}��>#�-D��Η�Ź��c)G��(]a?�m�+���y��-�B2����()W�XEx��
��B<��N�8�L���L����0�'Es�h�NX�Ѡ	��I��*�c�w�w@3��QA��G�=��	���	z�gk�_)�A���_�W���d��D>��An:P7��NӲ���\sY4ca	,��1�l���pB�qby����jn�ZK������Z���H������;�X$ߤ���0B��4��f�{�cuf��l,����$<-�m���֣��nkAm������v�N�3;�$����k�a���7ײ�hɱ���N�y��m�.o1Neմ�Í+�{a�#�|�����]�MNX\/�����Ya�l&ʹ'��ޠ���e:N�ܰ��x0֙���'Pa�����\۱n_(��J�Ԗ�ݫjo�5��4��֍���ɔ%ٗ��;��=�H�=q|x�D����&�������1�i�\9���@�4h{�}�ޘ�}$���o]���(h���)�p�Q/�ȞN/ߊ$�"U�k����(�m����\a���ʥuu=o$a�hCxDQ�=������^N\��W.bY�P�	�K���̥j���D��Y���x�b�C�����a�r�3����z�m��h�9����}a'���ȣ�&(�L�(�C7��������#t���Ym��/����l���ꚽ{Y
�\�*�?�%$�1N5e�d�~�S�����<_ҢF��5���r���H%�F����r���?���Q������Bncw�C;#���q�.C�b|-�`�Q׵N ���J��b��_�hI�^�X�J*y�Ğ��g�#K��>P���qUj�/b�e�v�m�8����Q��x�������m��Q��{�l2��h�v�-ve��o'���!A�.�������
�.IK0���27�P�83�bB�������n��p���e�R"�CDI�$T��!�j�A�׷�TM��&A~�����Q�&�f,@�0X���er� 4,8/��0>���¸�{��b��B���bFe��m�|��ȴEP�m�3�A6��m���K������N⃆ئuE�kn��R��c���h+���C릩�O��(���$��4|N���=����3f&���t���?5��e�����*~����F�1��z.��:�S��~�8�o�@8��0��E���mFK�5���)i�*�C�3B�()(w�̇�d�8��"��4z2�P9A�C�U'*�-���T,�>Y-N'X���'`�v��I�8q�m�ҕ���\w�����g���� ���NO$7|w푂F�(�3mg���l8�������8���̣�$j4P�|wh�@��N�Q�eq~3����G�;*��]˚�50;D���P�B��m>�PT{��G���>L�$�,?�9k��<q�L�-��t`��dN��' ݰ����^�R�c5�yݚ�Dt�R����b�J1S"�b�s��)w��_vR �/mI��xiJ0���(��
$�!wy�s�l��P56zK���-�QU������a���	bա��CQ�ɹ*�����G`����Pҩ�cu�K���D���sw�!� G-x`�(���ś����dg�Y���s˗7�F��Y���^��n�9�-b�T���ے@A"��>Dy.�G�2�����q��F��j�(�8�[s�o:�e=`��0
w��W~���I`�mښ:����u�)������,z4�Mw���Z?����oo��f8��!ߝ�Y_	*/K����wrp����N!��@ ~<�2D�y��3<��R�l��8έ
�{��lV_-��|�ò��9Ae̓��I�	��8�-��"�y�n�cH���L:���
3,�*���Bs�* ��y��	���,����el* �)�`F���\X��q]�՚��F��7��S�f�]>�'�'�z�7���z����d:Af'�4C����b��SQ�[�gȤ3\��B/�ܹ4�R�����v�����[�/�zw'b«�����dd�⋛P
Un�į�S^�B�� ���it^Q�>�&�0�@�?�E�z���!���[��/	�r�55����I�a@&����������������k�p|B��[}}!c��:�&��Ri[��aA�'�J�^Z!��ˏJ�W�#�c�.���L�"�9�!E�paX2e��q�;���N�0H,�,#x*"@Ìty�0%o�)gVe��j �ʲ8� p$M�in5�2�;v��ւ'Ůߊ6k�&҉�_(�!0}��s܉Q�]G#/p�$I�Ym��hxNED�܀iRVWB��Ȝ���;ásB��ê�^�\T�2<�9,�/p�{�>���dѣ����M���G'��%dx��^����D��s��M1t6�6K�!t��b���<p^T�7���(6�b�fٮ�ؘ��c�x�[�{����s��:U޳��?5�O\�����kJ�L��=N��%U^��~5f���_�P/�֙� 4*2�$SK���EN^&�M������[��_̡����ӏ)�y�`!ح��b��`�Om[�)aF6G�ې�\�G��H���s�Ί�"q��J
�-�E���+g;&�w�U�7�ڇp#�qK���	Ӝ�ȷ>"j��J�r����򬠅v�w���S��̉�Y�!���&~���{����;پ�/�0�z���|-w�\�S�磶gaMsR����xiF���~Ht4	��3���4 ���b���`���$�����̴"L��h�I�N`a���j�
�[���}���DT���!v�Yx#80҅]?t�m�����B�?�l��"mц�AD��C��t�TD��{���I��M���)}����-�۪�9Q.E�g��rt��w1�st�F��!�b	�r��:���j��[�O��M\[u�к?]��������?7h��I�,�l��T����uHن�E�����I�l[&g�����p�D&m�;g��XV6 "��f�>�Us΢`/�Zf*�_���g�h)�����JrIg��:����Gl�[�O�SW�x���\�$�yn~2��x��3��Ш�1Ԛ�{RZ����`�=����|,���O�=�0f�w���b��Ox�x��-��..Q�,�C�)����F�*+1����})��ѭ�5�}L�L�^���P�G`�O��ԉf�s�ow���X|�3��>�,���Kb���{p���ډ8���E)�n	s,�W��݈���ը�>����P�BT��IZ jF5��}7��\���5�x#�/�$�YH�6J��E>�%u��C�������)x�sO�Sʁr�Y:���:�>F��9s=q�'�� o�O��K-H[��"T�v���ڴ(����˽"2���v9Y�?Y��Xn<�W�w ]�#�����4���:�{MCѽ�n�?�^A��X���D.T�W2��_�)`rVL�V�����̺ ���v���$2����tADC.���>9an�%�C�M�'�`ث�B��Al���_�y�Q��w�U����-n�r���X�C�VI�.�B�k��פ��&s�R�	���꣇ۀhg��oT�����.-�6�CE�F_�u"ܲ�vɳpԦ�������gC
�'��1v�D� ��8[�ʻ�t'��)���Lo<�!�u��p�6�j0z+P���箤k���g���_�V�k�)Q�*1���SW`y+����Wc���M@��!�r40�s<��X�!p��n��\:3���/���ߐ�@�*T`�����a�o�ǟW(9R�9eB9E��j>D�(�w�t��vfa������������iL�z��Ӯ������U�[of|��Qe��|�Y���,A���]~c����8Y7����(Oo�=hM5U��p��~lN�6�BY�/e�dŊ'�b�px��	m_jo�F�2�;i�h�q��+�)���@�P�0H�zx����`:i�<��zPi�ӗ����q�hx&��%%fJ�W�R�J��>"��9c��ra70���h����/i7�8��bOTS{��͔T�XCvi*��t`.>&Z�2����RQ��v{�)G��~�$�|K����U׀K���e�6�b�e�:	�s����Bԭ*�F�A;?\Tem/��
�A�Ve�T�F�t��l/M��73�_&���<;y�7hV�Q��nS�y�_:����9�c�G�	7�t&���; �>�w�b��58���|�����.��(�،���;'�qѭ��5�ߌJ��0<�<vqG�&��`��c�)�̵��$��3`�hQ¢�MI�kR�N����a�h��K΂茟�c3q	BEP��#y�<����]0J�#�zyy^��t�<�lXd�Y��h�7��󘛭}���������@�{����v� ��+����0+�t~=�.�� ���9��}2�P��҈(,mZ���C`��1�s����9c�lB�k�v��d���[��`�%|��K�Hs5-����4�4 �@������ ;��3�/��U�>W R�Q��$�$��'H����u��ӈ]���֊���1g�0�8j���S+�&�	��W�8��ˢ���x��������I�<���!�1L������ƺ+si������E�����&\�$F�ߦ>A�'�"z�xÃ�A� 3�~��X�z�E�5��/�o�ܻKNh;�!���4q�QXX�p������?��uU";�����<�AN��@�[[�y��ٲ̄q���"��XL�� �Y����Ƞ�Ȁ�>�(��u��sh�ؘ��� u�6m����6���!��l�,�l��)�=u��k���*��R�P��㩽�� �%�8[�w�:�1�����C���rh����=�v�쇮~K��b������M�	�6��B�PKͳ:kc�݊ ����i��EZr�g�Q��p��r�.L+�A�/�]vK0Ĝ2�)|\������@����F��;�ry���|�)�6=��J&�c�v �s��%8:%~@��8eY����'�1��<�_�tTX��dI{K�rXC�q�M$i���҄��WtjFI���f&0
^�zY�6 S�_�a��4@��@���j�K>�2J���k+���O��P��<q)�u�29K���d�8�d�j��B�Qj����i�t�E�0�΢l�8�DM��`�N���׼7�v��{�6%ɱr�p���`4���M��H]0qF�? w1� ��8g�.ڣ"՞���w������zD��`��hIg~Ą�k���
�n?j�D�s�=�����ޓ~�k�4CT���#��
|F���8�}[֨����lU�Re�dg�0VM��ᡁa?�T4�3��v5�$�l~E������������(��	9Z����ǆ!�c�p�eu�{���A���$e�q��5�lr���J�vK����@�Wq� ���]���Az�i6�K�u$����8W�C�=i,�z��n�@/�5͆-p�+^H�1t+��Ԏ���%vV-�١2�l��A(���#�_g��6�y��/�(�C�G����ܰ�Γ����t�;��>{dU^��[@�ՏƮׅ��ԃt��cwr�-���Z�K���!+HW�4d4Z="S�7|3v�)%�h�sPm�ˠ�������{Yr�������jy��m>6�자���<CA��@��K��]�Ey�aO�ُ�v079�p��S*Ũ��GN!��(}�i	y�be�Ⓡ��k(G��j�6�WL��<̐U�*3�n:O;����Ⱥ�*�J�@^e��L1'V�(ȳ109�s� }Wm�p`D~M��R�1~0�X+�H>�#�G�����r�;���ʙ֔nŽ�8�*�PF'�=��\��+��e�,��̆E(��<&p� ܖ�{���܂TzK�� n�@�[��ز�c��9����J�S�!�ż�I/�;����]�oT�w.)5�_ml��DP.��2`x��d�넬S�K���?���]����i���6��+����7�m+QR��g���g>G<��ʿ�yE:T���lϱѵkr��cx���Ӕ����-�BqW��j�0�6�_jv�h/�?ͦ��>�j�t? a��h�g�**�f�Q�S��5�]��ˈB��i�")�⺜|C����Q�P�ha��&%5~�ad�U+ꆗ������tӈ]g!xIh;�^��8��I���Hw��t��F'�Ӛ�ÈZ��\L�.���s�W��(Q�$nG4Τm�P;ڡ%��������YTE����;�T�N��KL��E:
B<lq�v�
޽W�<��
�
?˰ܮ�5�{FЊе�b��� ��*��oց��Ѕ8L���ܭkY l��-SI���K�^a�H,�0���H�:��r���=o����������'����xx�Y��?F��?��@p_����Ե�()�3G�H	�4Đ�������fW޸�p��٩K�o�X�e�}�"���UM�֊�׬���H|��e��������b�޾��k;�^��[N��)5�f�i�[Ij�M�:�V$X�x? �I<� �<"�
�cp4A�C���\�s�`�K�H�,ʋ�>oW
ޑf��y����y�B|q����!����!f{�`y	�GgA#ƚ���f��;�e�������h����WMTߝj�K��y��7&JA+���f�sfI*k��m�|W��ϙq*�5ʄ�!-- 
�v�eQF�ͻ�����<�b%!�N��[���+��(����Z�Eڣi{�dԧ�
�K���N��fu=��ҁ�YsN�ɧGb:r���!���?�`A5o���1����4��=��lLjꔄ6�v��v�2Ii�O~!�<DD���cUC,)��%5H�����o"M��=w蔈�&�q{}�GL�c�F�;*��>���y t�-��:{F���8!��aOvb
C�#����쾃�u��ף�H;��N�L0J��?��!Ũ�с�R��a�sGG�$�	��N������!��Qut�O��N�ee0%����3j�Ɲ��� A�
�t��7�{u@7�#AFϳp��-��JT��*ҕ��PH�t�����2�@2%����EH8q`b
%��_���y���? �"p��ȡn����8Gv�j�e,���,Ua���_��6N8^O��y$T��N| Ë�8���@���Wd��{��_��-2U#"����i��FdB0xPL�k#���̶�+��vr��|�CIb[�ʚ�����A�����@���a�%��7С��h�ܣ++0�J�XX�ֻ��J�4
�����\,:��L)Q����$;
�!�Z�ʬ(\N�7����#���Or��)�� L�l���#	�ҕx�j��2
c�᠛��#�?W�%��ˑb��V�����qO����"*�{���s����maп�nbq�]��R*�Ǐ��[��0R��Ў˧���a=8ayT]tР7)#DF�B���ӽugb�%���|>wo~����W�V1������ʞ���������7�<�o(yY^7�����Q���%�II�,������f����"���j��bQ|J�}P�g��ndl	?�>J�E�e��ПjAT�i��WL����D/��$`ː���,%U��G����S�Y�keXƮ�u���� ��S�*�w}����z�Q���2�9v�^q�	G9N�֫�a��	h��������R�9�p��y�	z�� O�,aH�.�z��H�|��Ff���k�T\��:��Q���'ۙ�&���BR���bK���"Y