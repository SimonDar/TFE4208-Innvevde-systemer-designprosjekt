-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ba1abvPiUmKWubqjRR1u1Kb78m+GManOlwxG3onMbw30uijkDqdB8fC+EFEMcPn0MX90+mwvRS8L
FhVMtubM1yD+9vTrWXm+a45tmafDfl5cx59Ik+C8TvzLuG6ASf3PxaeUw0TrvYTaPUVAk54LvJN4
ideNfPjtKn7fQTEd1MH8klsHrXaZiph3phrKPPtpJ454O8k1O7PVqRLk4jaZfqmggWVLVzSEVfGU
uDKuFbsPa/ZAdSAdz8XYB0s5dn7wBgrU51MZTbEbeUUV3p6mb00+l53liScco9nS7jeES5tmI2VH
KMhRFZEbNQhSgRmACFg1cML0jYa4TUmaL3TiOQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
1DwshRT6SR4KUQC8KzK/GrtV7AX/Fw2McC5O/RUu/VL9CWWMx2WLkuXWkfUWPhzle4WqFr9+BrVM
L00P+W4lUqs6OF9tt8ypaj/eTAD1UU8M/AbdfgxYC8fD6b7+JS88zeis7F9dnzB0wvnxoeubdS9Y
Rt6mdPmlbF5TrkZ61SysJ52W+AidLNcdtoo6zDf8KBFrJuiX2h+0Hg3GyywLSdmUpJa8fZGorOKN
mniyy6bhS+tivte/IaTG/6nk2lcBIW/cGzQMjOoBk18jodPn6NWyeeo4Eb9jQV28/ZtIEdfJ/0pk
gPE9MyAw5I9q6fQy9m89G4/Wz9EWhHFPPYGKAXZolnf/j6Va7I/55lvHo7L8r+DcHYtfrq36iln3
94gffporE2g1087UUchblH4FOQv4pOgALH4HOv35BwVQyNnYuUEgkqyixxk2XI4tlf7adi1Cf8Xd
NJIiqG3NgzF7PPVCHA7NuDX6A4GIHLxDt275wnWhO9mK3TWNJ3HxqyS7E/PuMxYw0IKsc55vYw06
rhtcCDp6MaoUwgsRgouRhp4fgwQzaZdq7T6JZRfXkppwv/5QSdhkhNYV+zaImlrlzADNTskfuoXU
1J4GpafXsYniDUDEbJqFRvTLsPSUIK85tdlMdhwH/LyDPmpGMbXZtkzRCDipf4K2UKea98gl10Q5
Ol+7IKB4WKRo3ydaB/9SzWSY6yQUnADIN2SXiObp6bD6xo1AOcVRcPiCqOLBuTNlRbQwTDKtiG/6
VxC/yHRhwL9m7IpJKxxnuGBd050Pf43aGbb1Lo2QoBu7fY56RYJRNQLVhRz+ZqqHfM7OvcXDBPQM
TGsXvklFv+kmuQTzZW6n3tOWrhVmTEx1hePV2O/UWOJCBw+0+p+mk0w13VEL95/7Aa7iiBiKVmwm
GsaQ+pulYdZKbO9jrnLBUfa+J5y0uT7YhksELocTZ/C2hmwvmqoLgfNjTBaVkUCtkTz2M76OKpoZ
vay0HQAN73hHWn0nXoWHhaeUTtXtvbyuubkWK1WveUdzA5frTi0hH7JlO9I8deHc4zNAlsecPgbE
xCx7z9FW6Q7F9ogkHwXjqrS0OkO+K6Mi9zag+DQYT5no0GYOqNoudzT3deOXJRf7Jq4tqFasL295
IokYKcZybkSehyPD5/MFCEJFbh0I+Ztb6ErQ33twgkWn3I4Y4/2nJOI7fBdOw1clx0bpO0bKmgZF
0VFcEAeK3yGYGxZKkyRha8XkhVzyXwtgbfvRtqMDQthHoTJVuuRrOTxqmN/pIq4juQQegLPpxuOv
kDqvPS5SKZ+V5iOaVPNI7bOcBDLMZUmK75c8s6dO3beToshgAx04nhzK57UaASNH8bKn2gTwoTzX
W7rxFSZuQ+WF9lckfDFuazEw9Og3wOswn44nxCQ/2mkSAoaP65qrSYeIxmQm1F94BNgvctwju96/
mcn8XYyPCLPlpeTJyflz/dwSl64iWYillwGwLSeRj52YaW4cUpqw12gBenQj6aQIYFoKFkg9dfds
/JEUPVs9/k4pdyX/CsYNF6gjsnrJXT2fNFYrDs5HsFa8qv50okUqJCIc7xW+a6+yuHTEnTXlAUJA
FNJxyZPZL1Y4Q/qo1ynFZIuvAS3QZeTQBXiV7hCjz4omVsByWvVGBVOruMc20l/XwL0WT6/rP4Uc
Niu4AWd0Lcxllp7wOUgVQqhVzTZWJV7eR1bmDsWiC+2tkrcaK4wSSidYGnw2PX4nvbXXj5gAyCcM
z0+clgdzcO0V3JrObYJB5kDstTI30/FFlKPhqLE9PxBbQoJGK63ToMJTOIsq7od7VxGCa2TZgLC/
vc6cwGX69hWDghzaIgikzf80aanPHPxHDJL7xf2w4BJMs+n6srah+KUydf9B01LtXa5N/eVBqc8w
mojCYjmni02Xme+AsHu+A5JKjIyeNhQx0z9HX21OAdVjRaZIh6/9RfUzibaa8t5cP1y+BSoMUsOE
1yLXEfscwHcHEig3qk3xRUCzDlcPcAseXxd8J8Lwc/a/Tvn87Q+c/aeVvtzRakTODYzJ9kdNvuo8
YmKcKk8Ra7gCXN2HNGwQCxg+8f3GHSBk3IfmjS+bJaUuQJ32SDNNja+bTkMWaB09PN2fwUuLEp6e
aMC20YDuMaAO2a0SIPvhJTj0E1hxC54HJI2n4iLvz0oSSskfJQjLbAzoG2ZkocNKXNe0VfNU46ci
sEgJfycHe80JyMrzzcsJdc9Zui3P9tE2r/wjCjrwC931LDj/ThpsJGon+iUKa/qOzZ0C2HH0c+V6
muIaVXUKKpb0EKxHGloxOJj3
`protect end_protected
