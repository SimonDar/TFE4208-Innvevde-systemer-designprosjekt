-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
C5+jSJJUPcquoAC2ikUCItmAMiRIYKK4LzeoQttAS/p4hO7nkZPL/kRQrAzOqbPQ7+SVHixxsH21
ncke7ACvpSkgB3sEd9td3A1Dl15YcbyWihdhKME6eD0TI4PbTWBPlVZT9f66tvhiQaLnGSWi2mgt
CZrHlA7yGo4fsqtEOgxqEzJl1Qjdde9YLE9Vt8hZCFYHHKNbm88Q7B+H30UHHYnFL1SMckkOCVJ6
OcRxqNUJEajmtjMrDejMWeoX0DlXd7+gXO918Sv54Hnb23UddOvf+gBHNbkKm6p2vOMZbgFr0k8P
WSPRNH55isxFzCdKW8HaVUk+En44HtDNvw6/QQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
63FJ6X6t3GaFqSx4y9H5cjE/OqX5HA9hw2yw1jVbL7fxh33pxdczs2pWDSudx5skGkcJbMoEEHdn
FFI01Z4oNqzbyhpDtXgU9ClGDRVhMXZaKjnL9/jeYBjp+5rwNIUNxqN3AUFliWx0v/mc83PmylhZ
AySmfICcMWyXD1aMazHGGAmRsfgpLuBCU3dS+DhMuctYANPyqEsSl2Tm1o3xuZ1Gyn62CWvJWK6M
w7UbYMrerN0ksouwRtqN40GboFPxgEcyayzIirYm+unAL7glcXstb5tVvn7gpciFh1Cd/C8TWF2d
4dBiX5d71u9exjyo/nK3yFcV2ryDa+9HZA0V4l5N920hGCM3wlPe2cfOdHvA7iminPDaCPcntLGD
NQw+maMID5QHjnftdj8oL6OPXbROD9aPZ5OVvGjvy4pIY1bEwEdafab9Vw/1psGRbz7GZOOryUJB
87+uNypHPud5YrPzWYDzrP91FiIVKhZpnF0wA5XC5h6MoH44EOF3AXZUqGmLlPNNNPte+UXJbA6Y
leZrK1bgIKJz0DelWNp5+MaYqe6FCfhYzrm5yVxmj3H/Vdb7tcGx2uetedV+hyqH+jSoIxgRjsTn
by02O4/1LT7X5xiLxbalK6XzvM1QCdK7rnCE/tPgPchDE/x/LBcejTzCfeVMyPD3SQA8LLcxD12W
sSDd+stFUb6E9oyLee7AC/3u6JBsWDg27RIj10ST5e22S2eo1cqr1X8z55gV9jxJwu1OIbBNzHgQ
abK/ectjf/dwybnnNg2i321OIT4R/ZVDSt5yN29DGFy8sInwsGoFXe0kKs+yEc33Y6t0jB7+RjPs
3GpDXb2EeEJNH+CXPUi8DFitkQn+AUI1ogVIVNTqmcheoN/x8i4J2dqZNrMD7EZriGyKJhZG6Whs
ZwHwfV0ofiQ/Ex2ND7tMLR1B41m1E0QJ133WsIgwn+gk4AoE5z/kaTyJPOi3mRHLtF8ZKNeMAaRI
l6XegpYFMtOINyKzntn7TqhMXXD6vX5WaN+52nBPTzx68+LMyA3DtG1JYji2ywhNi6j5QeNR3VQf
XA8G85rzpMuaXizIyLFJz/WZqQw8zvEIfBWaV3F2AcN8WmTV32RLvRCNQLVEO1kNtibPLUguvHtd
DkhE/aUxEFw2MN+LC4An1xC/k9Zg3RftexTM/i/XRmwc4sHPxb9bvvQxk9Jlv+UKfJSW2FeVxsyt
vkFt37Hl0H2Y4gcoxV1+pqCc3arnOLiwBwaCiSeAQJD8mimjsUutQ1oKrqueOMAGjXdNUZ4entcB
530Lm3F09y8gVLR/xXgdNdOp3QUHRveJmz+RbXN7SiecCIkYlofsA7I7oLfeYjaE0tDdXrhEg+Ge
L/lz0zedBRW2LMsg4AOY67z+nqJZPx+rWUCDvS07X86aDNh7RXd8+XxJjhE0lwxBvfrw81I/OhUM
17gCTTfcmxuDCS8gsSWF4kYVr1wq1S3G1OiKwQslGea6Jx6G/0XJrJtL6YH68qs9wpvQo2Ac0xX+
4YECOXVEu4av6yQtbmNmrNa4ptT+cheMJ/2vOE3NJbi0BSALF56VQ8T+0NAb+5kgUvWX45aKDHRg
0u1sK4o8iNFYls7VSiRM+qbBHWllT3NYSTGZ7UjeaxEFEdKxR5jDO97jGFq1o2D09Xu7weFAFjul
4qsQF8hfgIO8wZGczrnfHKMmqaDKTRAIgr8Oa1CgoU4se+prIntU+h1VEUoQHfrifndT3EKHQGc+
3mr1vMFDzqFy7si9FAH6EavtZab17Vjey74Ee3hJ8Vlcnlb9gY6Tjzy3I4OyKaD8nhU+SSWOMAM3
8Ieh01T0Txc3J7o7HguBylOjWybYicskAyp8kBr/EDxyJqyReic+p0Dgm9dms9ejK4CS0eki0Zn0
65NdauetqoRUVH4NIqtjwNpY9gfxQxdyueI4CGy3E/Dt6q2QIOky90QIq/LjJb1UGh0hQ1X1zQ5M
r2GHpEgG78hlm//um1038a3G+DxbPGzGKLG8AFiqb8e0fNa3V9Yx6BgZ18YWcUCS9sABPaVuCHBw
VsPc630/PeqWBpOzE3U+P0lEogjJWvxv5PpQQbyjE/N1zCBuZz/4IqQNz93ACivgoh3hoErnFBQX
4QLMONLO0CMPoXwchQMgqIgTMr+S8/jBRRIhjGuSYBTkri0FT61I49ICpoDxwk7pcW0SbWfKr8R9
56vffPeB50ewc4iy0vKrMdIs/LeC3SiV4l0NNTNNch+TzKba80Y25s0GLN7bo2G0q/m87Up8CPny
O5VUR5abjGxeDPmq+GVV4c1JGbN7USFFY8n/GyoN2ISpvs5+g5a/Kk3B18uCGP66ZY7e+ZEYJRgi
O6I+S02OfFGWFCxS0GcJjr5RQqVauIUwyH47zjfRG+pJtZj6YqYI8l/jahCLnUkgiKt7AlqgFD9/
+9fNoMaIwdZWuldbTMu+lZZLuDxrKmmOvvNmEvCUCVIc9lh8q/lsT3onHVc5vK3DK/Xt5wLbGdDo
0RUXztdyplkXl5lZkCy2GyX4BFqEIieSRHKsFrVZl9bkR8ypEISx8i56oXNK6+dQM4EiqeeoqyK4
cpjjJBOm1uEszNLJbgpmT5EgDFD5LFzGJ2r0DUXvNOgIIlwEVNzbbMsVP3IK6gfjTpVhDbOlECaL
NHRG7gDafg/Cr3pzNugHLCvpc7/EstBW2oRrJwZ9XV65SNtPBOmE+puzuST9MNPaKIKChV9XUMfq
HTQ8uMUjVOkk1EvxfLT01tUZexIyYwSeBbefkXmw4ovvWew5JVWQsE/Z4TA3EYrSiH8FmeH2Y0HG
xzxOqBaA8aEA1Pz1MuFCa9HOpar86OVBHDs7AudTMlhu4yT7RbP5WTXDbLLfOTVrpFcGVWrUofNV
IEDxF73kMPOuZ18XqeUd27p4TSdzs70uwxEDWbUUEZljDzooN1Jaw9lW92x1iWWxGMzCoK5azlu7
bP49pOwe+tayLK/aPRQ+vI7rBAZUBp/4Q28nA67qZAf2AH64bHicFnRH2ft0sbB8jeUGpmuX7rFj
PeMksFjrnJ/N7y8C2tN3UCnimSvPrDJMszwvWwSx9CxYXtZaq8QGhYwkNOtfcMmdrmY/aT6OwIxK
ms7MKX4wUioloxCpOyeM2yAWoou9f2T5uTPwLIF13IcYChWkMegV8CXzATRlviUi2LAXJNt7g92u
t8gnruxKzzyj+atmsq7tyAkCoIzH/PniZMQrV2ZjPHlIWt6aUc9JNJp9XRQDhHpaq5nibOM9PSHf
f8WSYBA02c6DAVQmwY+yZ4QSriw5Jh94uJmH+PKCNp9xnVFHRX99eeDMi/1nM3fD8Lk6CGm05IbC
J7WCY0VIW6mqrWdmZlZ0yF2HcVsZ8v34viKlDlr9cyqv3A1hve0KFUxAHFCkLr/nRejVOMIB/XJ7
rAVAIUSPSEPXn3mTMFtlFEG2TvKZl2nbG9HIbsLbfWsx5yMQ7ffrYB/Rf09qwWOjxW2+5nZrLj5w
sKvC/U0CJAO6KksfmWsOOwjpLyE36Mtim6VkBmWiMSA0mMEcPcSQFbxGZxHduJJ2vyhzaO1VWEN7
zVA6hIT0zD3H1tFTs/B0+Kn9Jaz2gtTJ0bJZbewUccdNcAOMICG+rqjK1Y4RJan3iChkey6RDnTN
JclCghbVsqgfrxK95DFar2wCM/ATMc0g7fec/uKWMFMm38e402TeMZNezT7H92W5xbjokozpwRWT
iQvrGP8xAaNXt7aW2NHMisPTUOaC99CxLwkL5zvIL+1+mNov2HI0WQCAs5BLzNru4c49m5GOVFMX
zh36UrbabAauKd8QnNn0gEA3wFOVmZTXek7nx3H0gBOFCacKwEIBkYlGUpXlhLLP4lmac7rWNHFE
fXqB5ZeniEkrxYBpUqmemanMAdxaEr04dV8yo91Tu/wMltg1UR+kno6HvYEz/awdToFLvzOc/tmt
c3fPLAxo3dEdPyFBrS8F18ZuOH03DhDR9OFZujrZDTKi7QPyyQ2btYM6AxXnMVUtkE/L4Q4+aMUa
V7TK7cftmef3m8UFkmI2sRz75mR6n8uNsT+FWE1/14eTozeH4+2G72PL59LjVCItOWExYybP8zYA
icDUBg6SHLYt30AU3IGwx72xxQZsl8auowpaA/gylQnm1Be5XtpOV/y9Jg8+dYPyrCuUcQCBTxX4
zKzYfZc4uGxzjwfi2fAYcnDw5y/6+M1SToohI3I86ulfq6atwFXJ7AUml3KnbwfPItwDXBO4GEmd
wv61ikGlRFb8dZH7FTa2Dj+WQnyaiMFGYgZvZMsH4MVOz/iwDhZ9xjPUtu7KUic4IENpJNv0f6fY
Ua8/iBF3YA16m9Pp+qwMI5VaKCsz2gO3UcIMpRJEDCZ0WXPwAByutIBN1jK1JnMpg3WYnx9RQ+sF
9hjT/xVS09wiMBHUwwUjBiElaeFhFqbYabWGURsP4CIYffckBIzZGibKye5xIoImCxO9thCr9F3Q
Y3PXpE2hFEKvzv5FdOlrATO+wEAiH7TIi8502BGDJ4cOTiaxuPB6pWqmqjn8JFeUhWWSTxOnPdYN
ZbhuWpV2pumntElbDUHTlf2xvdsrRCeOKL2t0RVgmXNfoBCLDqudLueSI92Moal+gLBHJvSn1a+J
W4DL5NybHl2H2lOc6gpyaLDsoqdCxXYl9lg7MA/tfogn+ulMGOg16yGaz0svTMDcb7X8k0jsGdUX
h09Ffp1f0M73Vv7NRNmTy+ylI1BrHVJMVw0kX+y2aiu0SE1P4G+TykPTsEWE+ltC8ieO/pDuEb4w
mEascfxuvD6wcaywTaawOh5/rtCRU98DIoAOD0lCQnRECJKiCPpNeePmKEKTZriMrB3cd4xm9KXR
SBfowBI3Ku4vw4jB+ueyifvMrpWHqCL1Trfdu/pbas9x0b9cqLT7Qvx1RtTfKg3BqaSU5lQa4das
Bzw/VHAx5FZ2cxMKThKXZMjz6GkXLLW5PHt/yV2r2SoD0imRP1DAXtVEBcOvXCa6pCxIpMPQBq8l
v6D1jIWaGfhmmWfjEnuyUKjhRbfzXlka2e70ybmWzWyZop0DVtE/gcEmQ0DRBGFJ3TaVmPBiARWU
TH3XeWDNGJSGZdARSijI/4uvTv30pORMeg0FfeKPcnYmZT3BM+igCM+QZqLoJi16K5agiyesqLBr
SqluBCYmxw4HlNuyVLKQu6GQDgiBia2RkhAUnoPDMMJ/0nrHPwaJ0kMV4pKZse0NnvukmA8MTg/T
OxGz4ihsyFvB9GTFl7wOhTr36rLq0vd0mvQCxNcy9KOp8H8vaXmndr1yK7wbcwvFBzswblfKEzRJ
PFgljifkm0GLLmG89rfBsOK4fga6X7fLfhXybXWziOkORR8d0BE/Ky5+uHxq/mFKx1BisI5NToCI
XmiZZmdZ5/aHZA0oyr+xylcMgW5I1aQWkub7VcUz9roIGLZ0hkGU6qG0DrKnOE+Cf0HqK9UECG6X
1O8l1qXWjd5e50imWL7iQ40J1q62OEzt92A5FpqsbRipgXsu+k7oyKm9S53y7N9upGLv6SunNTcf
G1U1NSPZDJae9dFKFJzMegekvHsgevgn8M3U5aRbG4vwMGT6tMP9U3xp3FIWDdOgj+3DBpVXe27n
ZzxOld/UyQI6RAqgoTAwh27oScUQkzGskNqEIrhu1r4eol1E8Lw4PQEVuVr0cstrANlX9LqJJKZW
ThZ9zPjuD/qGaPzoEkN0V3cj7IytrHfjomlmhKKR+H3NNbiimEcrVRWNjGo9BFYYfVQZoigHlYGn
CnA55+1uumxXuWMz5p8qwZw8naS5NUCs6BFby6QNCUXQ8iG7gsLy05vJbMm96EpUrnzs2pUdsc++
J6ESqj7TYTCu5oypHM4l7aHfWm6jDRnGFK/rVRlyyhx9W6qKNWQEUtXJzz2yOmv2R1l2IDMjI873
j8GY7mzebP2vOnqJ1Mx4DIbxHoyZgCY5rTDmQYLlxwzYMP5FPpWDVyNkR0Qleshkr5izlLD7WOaA
9/D6Pwli8sOweUjJDQ60FLStPQADwcI3x9BPMXgShrjSQpWYE5KZY6qUYD6+tDektWXI8hqgV/NW
eCY/ZjQjOGK5SPIrGLEHutR6mVzBJSPGD/ayKBXIBB160Zb+fLe1aHQEuEjgaqwdlhdqpVXqZTFo
cwlThjpuaWFjVE+dOdEYdvY5386knqNv8Irt85GpKpBMzw+b89zkNAEw7qG25Gk3CqT8OdH0hoA8
Yb98KV4Ymr27Ch7rVfQwVRpgLnHEVVKOEkXvAKAkcvKKKrYbK4oByRKD6oaNPYvIidAucFJsp8ve
KLsPCv4I1id5SIImm2wrySORBhV4ERUu6s2iCI4s+5b9sylZD/jYJ4rYB9H4K75lfAfC51e6uHct
S4ggcUPoLzLm+MnpILWt7hfFQY4Rai19Jw0MfByGM8pIlHlAEbiejvAZqqTIvLM4LT2zYXn1QVu8
br9b1Tl4pMrKUXGnQtfwG4XC9sqGUOdrepzhQykp6AS5Ki+Ig3vLBOr5Nu0zqesOKx6vM2TDOnTw
yb0AV9iDVXl8FB4WMCPiCI0l9BO+TL758vRJBlAZ6cvf1pnlUGYZFlKj+2DueAIVgx9NlPB+1EK5
GgLmNRbbK/QVxwSOwlSMTGNqYgFSfpSDFojLSsoPEVma6ookIWzcgmFk6FkoeVpiUxXRNDRbZpHe
2IdTbVt9vbvZuSdeaHZaDtQybeK1TXZEfpLe232HOwKRLW0uQ43ZgDp4wxoOsoABPxM0/cDddbsd
R7Q1Ud3WeI69zu0JsH98GAprnQcEW5xy+TnUmsF+Ml/aGOgu3SlIV2NLz72fFX0lycFtvVDoHSO/
mAK+4kzScGltEyzfcSiUjSlmHv3rh/veNxA4KnNOKaloyeB0qfnM1b9aDV4RLelvu0/NaP0XQJYI
4SB89VS4PiFvTdjl4q1nhqv3iC1U08ybDwJYYwBOLn/zI3EAWxLwZ6rDXicbFtwUO5LluQK0cN/P
AjGnB86ADC/tT2gCMrwIUFznNb3Zzr/nMt6bwK4byfntPXN4XKHzD/iOAbBGWVlp837r6AAnjARX
sXfB9CxuHiGz52lAJEvmnNwohSYOAiGSDYDwkJDYmueb097nU+ZBpiV6Asy/9QohThYcGqihhkrK
gnNcdOMAVISzZZtOnv1qY/0a7pipnXCALF2knv0YephkzqRTi/fILm1Xp1hehqUwfRU5KkbsJMps
5Adh/8wIZbSX4HRex1h10sHOXAVmvOSdGnSVX7IaZZn4MrklM1mx6O+CtKbLhTWoM9klHPQYIbWW
GeYja66AWQIbDFe5FakdBlvP7XZ8NKe8ekePbeVfu5dTM1wRTI20Y599vatmA1XrBTRS2nmu3gAk
Vjf/ZB/J9+WgkmRFuQPwWvHE3rpdCA+o6jXN5dxEEPJ6qwPcFqiRKQ4vXu7MSTjP7Bvlo3xav8m+
sMWd/K2PQKabrFkJj0c3zpUZwokQKcvPoBr7YXzZO9KonGrgIZ/RxTi72tLkyLjUhqgfH8AL45XC
X/urJiiG6n1AE8jfENhsY90/o7BhjJc9EmRyIUYDEvUqdX1YnhLQXpueUEDFGXHw7dmEQD5WtOEK
pCM3F8ayXJh7gNpWrVheog1AsvdY9uPGPECaaqG+mieS5EE1UM22hRMFYWVUiCcjgyvAPTj75JqI
nZn27QvACB2z6GREs/MN6LNduMwNmx78+ORyG+Si51TYNT08LPCG/CHnPGUOiFvc/3UtgKNqSYP8
GsDnGfe2RGAlmDI7NJw4T6g56jlmctawyaDTyoVeADr0ShdzkOXU1yJb2IxsB9CKT4mK0hlTB+JO
1nkKTbXWftGbrNuyXs0o1WhDwYf+/xefomj4WWX6OiE2A1NoyYr3jswEz0C7vgr67ERHXoc5eZgW
BCrGee7mRNbFImLZaAgh0xaqpsG6YZTc1+k4YXJeKRaeZnOJk6eu5M5aCjBzwPVmfGT2ebWSn+2/
AuOHs7nqyV035obZ0CARGZPlFSZuut8Rn73j9GYvaKVUBJL0wWARiTwIdjW9pWJaXcUBjhJtRe/y
fckYDdtPqZBoIzBgwk7qczERgp9Ek5MMpwHZRtGSw+WuxnVMuKRViE9TBrhkqeWgY1zpheIoeO1w
EetglfA2DywodSU64AHRw5PkGr6jJMynMfackHyX9d6kWnbe2+7I0XmCf1Sb9pcWtrAD6SSqE7y0
UQvaTeKqdO5ahBxBaZUjS5yy5FHEDnYO5JHL9YLyFBhEH8aS1n0EsH3aQyCBDUx+ZkuvY8mJZ/j4
Iev+kaMV/4qtvLFFUZCkhcBfrp+CRAb/L/c+V/pdOb9shkToyKdycmpQiin4sXf2W7eAGiOsKtRC
rHZK0vX/Wa8neLO3DIlsZEKNSA9IZ4zmHpZDNjaOFFC9fy3Pr/Gs1i7dlnv3GPBSBtY48UNCb4eP
UsVZdvbp78V4TT1BgpI4Y1zn2wIonGm1FfmT+4lSeX2W6c3Om3CQZqiOVbWmvMGa0m5FE4oYDgM2
EqMJSNINah0+wRl43qJ8AqQ6SfWmsVPbj9GyHEBtXxuU2byDxVlYmnJQK1r8Xmsgs7ocRaZyWmOa
MIjg+QtRS5AE0wW6IG83XA1neeN5ZJObsGpY9Qk3HwaIis7UiRIZD6lgtPgOOw4tmevbK0+G1Yu5
VrFO4gN1Bnzl6w8ZPJ05Uck8fI2SJ+GypPImvMpmhFaDIy1ZOFTHCrUIC5vcU72DIECN5pjC/gfZ
NHGZkFaZxajS4nIrKvf/MwPuR0m/V5IbQvyYkoKKOfkTUc3BcW/+ewfquqplXoTq3wrRn0dxULQh
vPMxWfpZ1kKfqUL/Z94PraasperA5fxzevSmNsuRG/oSnKbQud77ZjmOWhYj5E9vHpjyQICbhQKl
7qo838N7nkCBEWhKJXPOOALDDt6HIlrTJou1xY1EiNUXDGc4gXyx82+flE4JkoRxwy0INQzc7w1d
qk7Sb1UMkkMHi4cLG/Jt/vzYO/Txbzqh66DF/tGV+v28Ln8D3S5s20PWujsKMlNWlhPtsOaNQX52
nOCqCDYyHqkpTAhsUkdx/+EkCzM2mZ8MgtM2hZktigTXWlt9fUFShyvC+rdXYq8eHpAUbwGsagMW
n9+kxSrMnHBmch5/ZRHd70m6PQTHqWVN2Wa04iSElij9/IZqMBk7Q5ffWTuv7LSMm39SsaxhfETQ
9U7CnvnUD2xfPh3V5dEZFepKrml981KX43fS0dPm8BL0dhisk1mwx9es6zNp1BsKrzsvJc/GH4IF
NZGz8EGcgq2aob98YhimhPKSRPLzJGFpOIvFJd2t7Xu/tpnLNnrdX2vLIG7MDad2dvRdLHQ3hmgr
vmNy2GkBk1mVK4nXR4OR3QkJ6Mh08XHjrKTbiYZQksdWeTacyihkUbnCJMrYNqSax+ijmQ6FYE1d
2qeoCxIQ/kCwajTrEgGvAqbwClFtLnUcA8FksnZZ1XncfkWOtTK1MeTKULqTZtoek5aKAlx818Nl
IPby35s+/1lgm3azK5AUt43dsets5SnOQiU9QRKXzFxDHMs10S8tMWiBmZdWtPwkc1SaELDXwPsm
aRn2XPm2k4KxhBa+UNn+vZW8YKdo344veXUJ88D8+XDjPERLhcH1skrRXUgz1WQVZqO5+cg0n9qZ
n6URUhV16Rmc5TCdXr8eY8UgL9kbaaEuEdTLytdHt8BL6RF8SxTQnklzyRXHKeXvHfLVeFA/ukdi
wKPevpejRmaujPVovX5XM5TwgzOymw+gKDSE88+fQvocHtIxvoHZfGc7Vcx3w0u3x4uBeMTbeJll
XRJe/NWOecwLcJKGy8jQqbjrRLYkjcxA+7SJV8YvIJrGNzsBoXaFBcVV1xMfxEYg0OK7NJP53JxZ
bgEkTwO9xJPGCdy03ANdHndF9pXthd/UxauPR8vKyz7D+ZVUZeUY0l+PY6TtEnie7qTSR/8ak3rl
AmT/7N722FInhahRkx603Dhs5MAXYFZwQ2OibQMHsfVjaTTmsDUsH3nv+jgxzOqMNwUqew/SuSgJ
rTgjCd5iTWzvi+/KqfZgZnKTtRV4u7ewIGv4QqcuHLNcZzNm2MyP12l63l+bNZTt0hi8GH35955g
Q/xS1Ia4YVn2OSlUnyP3mBdInPNch0XRPh/dmR1ihdUy5Yk0OqG/GPpgirjFvLjc/g1KkB5sSJuE
HYyZqKvzhHvIiu1cvYSaTS2SPkrlcZuQyq6ms4yjq+fG4QvFxqqa2ydBh/JoDN+YFC8BJoGpOc9c
jg9bNOlTGrxJUYpARPXjCD7S0bAt6PKpjZPwl2DLCkfmgAg/FJhYVNRVKB0VPslQlNYujqHoWuhV
K7MUTKlulKOwK9Ho63M4x5EO7s8cgetOLSz3H/Z8GCy6QzgU+U05sJjLf/JDU08RWOE/1gabiprk
boY0/eVjUg3i8vN4fDmBFrevKWCRLd+fRy8UGnNEDhzVqNimsZKUbpVO1QGttflzkO7S6Oa73Aw9
cbNXSJ/P2oQYYuHYQUt2lpNNuZtwzdy2tTjbauigRYzfhRMBFq0VK1xsvhZCRXLH8v2qksv6PAiN
rOv6MLoLr/hJxm7EMW1lgCFOSE3g7nExrHOdMhhMQpPhKvL1Oj9vXaAIWYV83ibfffk8ZDv+9e9q
gctPR7JQyr23Yk8HkKwAs76n6SIlqAr9Iglw857juiGfjwz3zwT8s2wNBxSvuiqPkHj8IKEuGBfO
OuTpZT+4/EtfWacK2WP21WD4mCzkwEqOKH7xtnv/kVpgG4gYnlaS49tvqQ8t8UGlaYYQMdJu5Bwq
SGIP6Ovqf/hzjcKuE1PAcm/if2FSvEDvtc95j3mW9I8woXCxYWau7ysw28yL1w3Oot3Qwnu4O1bw
JnZ8I3pxRDZwJ0BX9YrasznAJbKcLu4V1GuuSkkHyVfGzScYhEpyqQabOOtHYffxx8MJnWkAv/PU
sK/VuwFf0X3P/P22kpUvbMqTsbNaqu2ZYhgNKJes02vyGRmI5U7gYZnRfANjMoFwlb2uIBdSlCzm
kxoaQuBFXOlQid+L5TO44501fHkklViiKwGPrX66EVykDgBlLuQKPAeHx+XyP334EeoOZZcxNH5K
8BGMo2NOlp07RUQxzir8SBF13J3TwZq9D50B99fLNQw025MrHkok5Hd2e1DeVl6s7A01bigeMrF+
jNDUpWK/QadBF6Np7fiVFdc0fxIKGWt12qztp2/jtKcGzyTozkgppuA5vJ6w7vsgDX9dEZSiW7P6
cgAPVAJLUKpaf5/oeROKyJfLH4xrIAOOyl7buXWVz6MYvnG2KGZ935K8XzkjxmkEhDNKPvDhSaUu
FWwymDcUGl+L77cCZSksJOQfnSAoyKWRQGqF8iRoA4zOxbN3QipunJCN+8IL9o/O9HwdatLycHnY
MwXnQbR1Y5KxU7t51z+6zA/T97MxLxiugg7/btSFAdIny4fzZnnVT1q/7sFQDvqochOWYACsEUHJ
pwGwHHa5cZuqpYI+c4Y8PUI2O47D8YpzSfYCsQSDbXpeik/L/BHMpY26Owqwm84mq8Xhg2AK5AyO
BhIFHJ/Ksgf9BIS5b3b6NhIZyHmD9p0ylbdkhIzbvrPdua2x495TCcxU8kQGnc+H0KWBI2wDaPJA
Okkcvl1J4AX46aUw//m+TTgtuCnpj5gyMVJUbb0smQEk2588BGFjbRrwd711WlWw03k/HvgcRZn8
li2QqTxv6jydPM6eE6rjP8erz6q3uYkBk1mWANZcYTYsYPwEFUsaiXzxAy/4OUAuz/HOb7t0ITlp
0ncaHDPUPvTgw7hVVgQznC7iljF1+L8XLd9B140Wmn08QAaAC/UHWdwvYA7rMD4ukcLct0arOOzm
TAY+j3PhffTEvTIGExfmvY38o2D/Pqirji/rudSVvKcr9wgfWsm7gREZPN425wUKyoL69uRNKYG4
bMlbXzB11V9AZKmRqH+KnU3gM9rq6+Zrctjo3Gvz2acedyVtCCa4W82G9kUz1S/318V2smfZr7AA
ru7QSFfnEDdQ5Ebfzj8PhAACK1ttKl4J0GomwC46b6q03gkhlsVKCOWIHdMZhoo92BpUH78Xcy1D
uhS6tK/EPfnzzpZ4V4EHeO9iDj4RUK2PHZ/Q7iUAWfLf0vS+rqm06ik77I5i9c5RfJARkaNwrk5e
6G1njyeAWVNPePvrZs3HlGUfKK3QshCIRdYXMx0TUI0IadISxhzhiKkqhdIEQ4wEyVd9n6bIOcyx
kf7EgAU/spU+OeDp2FR52M4fFnbGb1L7p+8ouG35iO2s3jAdGrYb4UcFZhQijhaImNHG6eUKRGOj
AbDadufvDDVJTlV35JCYv0Z0ygbM6K59/ebX5p9DcvNalBD1vKNup/A2LLyc2FHyWqa/TrOdwKwU
Cx9VcnPjlpfC1FvFFe/keOmxGGpiBHMNe0+Fy2mNTbS2ujJf9DZI82MILrIIvA6lf5JXmthXFIEF
fB8v10Aw16eFaHg81qwYKUc68Dk90QauxB7qovpfwQt7zEwLMi/TMYw05qajO4Qv+HAS7f45uwwd
RVkSGvL2U6O4qth9U1VQGACQWmZ4lR1qJ9x0nRviPaSJNuyYI7D172d/a8O7/bgLwlSpWVs0Wo72
pwa8kRH+KHKHzdI+t7gYjToItLhUtUhRZgYwlQoM4LXAWbBr/UcxsNZNiGBVwhfrDt37CP+RHKlD
DhEPMw4hCju9e0Y/sbwg5qFRREiD8qiu0vQmmsM1uHMRy9uPcRmBMi1wnTO68PN/QUAQPHnj5yJC
vAlm7mxsy+h24M4uMpFL6J3xJ9QI/uBMCVRYhglFbjxPqv62XAOnk2vO5rc5GSmEOpMxEtduAoxo
OjKfZ9gGrHe31KaNp0SRGzY5qh6liaMPYauyjY1Oz5sBDXjDn/avqrn11aQiuzoBC83YgzbzOtOV
GuYm9v0MJQqFSeN1763EtqzD45ioR/sZ7uK3jYvxW7j9T5zog4z08Qkb5ouu3K5fM57lIEa/3g1E
u/6vOM1aPV84UVtQku3GkuqRqm13iCOw2VBEv93Ny0+NFHihXKjiHE6Up3m04ZG7NScI3F+73b2l
N0g6I7gCo9iKlSt714xFoH5RRLph7947qfVx7ZldjyLQFqucxh17aXZ/w08xj5gMSjTAob5BKHeT
XsF21HrWo3MW7v4fmJYgNUlz15kHqZJBuQCqryek/76LLWFjY4qMU1cey5R28DAWD01huQfi+9RF
HXtoiBB6e56laCbb5GGa2xjQiO9mLhlLHicEeRqlRd1wAoa3qBhtZTr+vzgucrGRwDxJ2gwnBsRC
H+pwFsD6Q1Uv2+tVXOH5jonK486kcMEjoKnZxW/CT7/ytMYNKellQL6/atGQH+qsIMPKD/LtD8LW
hDI/9PC9UVX8WOR4la5+ssJ8KRqZV3ahCHQ9cQihgMT87tvlTiyejDVJubWVCw1wB+PsTdkuyu0z
WLrzkVOcf8WdhdYhI/1PUa0GhwtKi5eO/MDq/IdqTPQm1Ennd6sWNp61NAt0QU1/5f36NUYSsRsT
KvsflFs3mU+LnmMZsgocNXwGQnjWMWAoqwb9fk0wo1gXrhtuXdGuwPbIohcVKLgXKidvfDHBj96Y
htwQmKLQayi8ngd8IPmkgA7JiZjDoU6ptPsIqtBk0Dz25eL+j0edSGE8kvdnHMJTzaiVGiD0d8fe
tm8gwfC7alSyWHdGO1EDuOt6CDYFz4fpTdW2RlaPkkCZbDcBwto++3huhlyghUrlaNSkfklbLJ1E
0SN7Na5H3exxlbBGnrQn7vXghOpSBHW2rEi7Y2P/OONofM/zFyRSC6QGHYqFeMdUPqbRkOw2j1fw
OjPBSfReCy72eX+TKidhddL8CpBOGTawDWGuLD9igF4t0kJr4vJCBxcUU39inInYUX1TCuyyff9q
k+rXPBb5DAWQGeK4DXBhsaCzmk9TnVLo8nrqsNKP3sGBcC656HuC9liQMVAjlQ+aW3ly354N0UBV
GBN43JwIb76AVLuEgbAtC4kA6wAleWJ5cbSyzqwS+8fWcbdYxUDVdndMmPVG5mIcmrgEHIRmWzgd
7cTJdgXe8EuFgOfCLOkiWWhD9j5JidyL6Oxs1QfwaiNwnM5VFp7KTJHG/VgOxYp9amXtDP4WvjKc
MVnLZkaX/KUS4mWGwAXIXyeq4NmbfbKCsx+YVvJaH4DHOb4Uw3xBpMA7y8/uCVecmmK3aaC2B5aa
4Jd+zDrEKxQTp7G+bMFs2N4jO9GUeGSJkqksTyI8OKrC5opX+yR+6ZaVol4p0YdSprIgRJKZtYX2
YFVtSE48B/TJxne28lc4120zol59hYJ+E6wGbHvfWmj37F/mlXqv6cDnBTnuWeWvrweeCGx9c3Zb
h4xudIkolyuVZnDsKDDogAe3qdVsT45rPa6APuM5idY3YzUOQxWVdtFIbcXgj4UEq7+A3mOqzRJy
xZcutLsrrDmeCpHwzVXk7pZZNuI3bCEEZB+RMqXrnrhf4SE1IB9E+86S3Q2euHbFOxnhJ7/gFoLD
GKfAPzUnckvCyjf4yXELk7qaYfcveYTYotvkN+dqkqKxpeQVlHETWNNeeYZ7DQd4qGTR/g/oRwlJ
3jS2jloqe9XmS1uDZO/h6nRUcONh6A0JoMQEQeWvIAbn9CHalTFKLQcGB8hRV8bDcP71EI2e+d3l
4jT+atqEVS1Oawk9yJaQzl/e4bahaTYGxcXA+9UM8xH8QlccZ/gep0xbkyPLf0YFQrIaXr+M62YU
8AW3LFQ15O1gTV3mTIHsNWiCio8pGo7LmUceh+UOxeQJa0SjeJKeXAw0n6GLSzbUN/5V033WdAJj
IhrD6I2qiGxWuHQGaiEu+1Q10rGw4Dm+TG+WnegRLbwd9kvWguuMiKBKirkZBPh0Z05m9xZsimVl
kJV1kNxkfcPUTpqKA+wnkfeLmw6wjqEsj0UjvI+MBwwh9+ldYEryZlWzZzuurTy5I1+PZGvy8Frx
CnJ3Cm+1ErXfJLhM0Qu5d1CasMKKQzQJbVfRJJZZ8GF8DwTryKfC7CtcIfns38MODjCneYlq2FKU
DMatg9rVwAMuwa7DyBdQOXsPHjins2CU//Fi1lIjjOVU8SkrsWjTyjjimXplp9iRcES2O27ctY5A
5o593OyrVV8QouNztbltUXyuWNzb2RBAT1VSFXbfBogeRdiHshzq2RdLTXN9y2mSm7R6bChUiMtH
fjdKLukDEbuIeXjIhBx3A4rV2DElWAYIxNDEvu0RZBgHu2q193/WhNnL8IYZy+5uDPVMwaBdlzWW
V2Qmc1GGeIuLLjEMBc0FEvpsroU62M4uVUz/3bNMIcFTELlj+6Gfl6m6r20V+EU4aHmtPiEnWBW3
+tVhaXtRhN49pm389ARXAAmwlpP4kMRlppqz85TK38Imiyfgja6/cF14OzWZCWEKZyj3/wMzoZGt
JolcNeGCt+tjAmYyRAJKNdu62Tz9E7y4wlPEE7W3hFqmfeW+5Tl8hYpQdWUdpu9Hkn04cZ/80YXP
8UlEsA2gf9X8tV6vFnLweUtGbwYKuPg+shrnNf+WVNPxY07Nkm5xRDuzgZXErNpnJ5RUeoNYR7SZ
arP88MVVbbUqSJL8qV30LeQmwA9vuLGnzinWOEQMvvPWdcNbBYC9Cvy2IhGB+dZHjyx0QPZaBpAN
gQEy5aAEMUlvPAL8wfgaiP/AZXtx1lk6N8I3+XVwY2SDKbsFMZoKWg1N+G7+vab3gerBg4IgM18c
kYrhrgEpsSsieIKacuzjC3BmHid+YLyK7cLOaZRBXd4+GeSDmrN5DzMVkSndix8zmsj8MB7k0yRt
7n4fFBKyWR6QRe2aArTwO9i4WpRd1GoSt/EFCTkq9QyYG1LtrZuB9sMuNFFcSE36BCNHrmxIoDgx
Lxyksq5lo70j23IV9PwBpJaoL1v4hr6PJFZXFWA1rOajJsYpqGeOEPkSzn8Q0oTZtxaERaokGPy0
2YuBdUbaWGRbIztYFCZZRw4vtlxLhv9WpLf8UC6HETvtl7GFtc3Gzarwb5j0VlAd5fungaZy9W3r
9ecaztSLnxyWHIMyU2R/dLus5UQ995cVj19zFjYp6ylRrBc3LXZh+fCgsmBcd+SiJ6XDEpTJs7Ak
ZOf08Lr/G3iMt/39yv3Q3h33fNz6nvD4yF5KsmYVgeif0hoI067R73Xo70cG2tp+o2FUT0SMnl/O
TYWSVfX0nSs6BydRkZTYoMB+f3igJ/MUXFvtHEHAWR6HP2ZM3cVmAyN+d8/gZxAZzN4zJ0Dl0U/J
GBz4MmBxTT/+BY5Rd9iETwbetgzMOcap8NG2lDZH9gUKXy+NqArKmW/g86Jk6fjXCRpP6YKuxx3R
4zBJfa+16bQv4X0R9pSAOavOi5dS/fx0UaD4eO9d25sT6caE91ea0tNweXInbmNEkYE8rMh3yHsE
4C/vUxc2etjMpaAEknPHSDMId8caCbs8q8yDEaOtN62ykhKnJd9PAR3Gc42xh0T5+ef50ybNqNHX
2JKH31awy3Dz2JFwXYMmH0A8YBtv59dkR/yWCIzfwWyhefHdyIZ8FlEVAauTatifXLjA/RARTSDT
LEOen1ZNoi3ijg54eBDlHfoW1EzUeE78lBKSvRae26XOiwv2D8vbd4cbASxx9FzP6QIFtYzdWoJd
vyZU3sVisY2LLsmeW7a0DFHa52RfkZotpOAG4I8kSpr5/iUDqmvXFROUjn0VTxSiUXonP1Nxxv85
NFYOI6GpLZ20hdIFTLW8bQJh/1jIq5awyFC2S2BFf4aRf+wNIU/RbORbCtJeJs8kRXAS+iqW0tHM
nLZE4ZwvdRwKy0JUcdkGiiCu+c0RB1xzsnAeZ+URDNxhDWCJhPVE0C7wHxrOCUGKCnkANWT65NJb
ra/Sxs1Taecb9FC1BqLpzoeo2BmIz8v93tP4reuuQhSgAWxFECE0d4NeiMqeuO9SQaTCzVO7XtqW
ntWTmKEnGOURxy+5qsWdXzWMTbviqLCajtL76zLcuGTnE3oQib7uSvajbt9qyEhytNYTEXyoS+bz
YCgcVlxHLaQ1tixRV6uRLdk40Rkv3/RiU/UxKdnOr3ZeoAfm3Xbe5ga0HGHJk7TsQAXc+XKAGHUx
5o44BJq4lAVu/XaR65/lvLIMmm+swKro+bay6bcoIeGu1buZCMdSgglQW+GKsNBMg92uNo+ZzCSm
HX9DeYeSmd0w1eu6Ej7gXFik1OOUpfwp9U379U8QlD/gxa/9ZXBZgIqWA479RqOUR9LZfxTh1XUP
Rqgmnc9t85DuNaoLuKpHdnUqftcczt6MMgoNIHQCj8iB9aGoIR04lth2PUEefWZvOdpzQnYEcOfP
4hR359mmj+OUB6vI6Xzvp0uA2AmsFkab59aHd4uN3mBRX/2e04tLSa8hTvlJdl6EcykzqigQnEBs
ApehRDbRjPc1WRGMkSZdhSDk6bNozrdJH0/8v289hRsMxRGNS/Xks2uAGDUrzw3sB3tICougnYFE
azxDPjWbKYpzOEXXTEDg+5x6sVN9BAaPdpmghKxRrRZcstH2VT+VOoi+w+oU6h9POOgfKRO7pKt9
8pzLRNqASxiETwUmli8/nBlYN2Ca/gJEKQVPm5LnsVHv0yLYh1T2vmPXz7EQCMv2Ao//+UXzoCeI
/NJXTe6JCFecHxPoK7rXDUNkkjit0oPJvpQp47cXLHWLNv+Scw7qwHM68bgmGwzyXuF+0K9i9Mrp
oAt6GDRPdepwRKWZVomEEP7P6eTKW6SYIijXFoHgDxGPOLU0yIAqMwODpsBcO3ETTGV8fO9eXA2w
9AmCaXhGq6ByLp5ovjMA2HHUOOpyU9pO7+QL5Szdx65TGNdnwcSxmZBdUqifxSYCcjb4FiiFxQX9
A2xVjmVOI0NXlzMZFh68IvzVpncaDlEsYpBWLOAyG/2LROw+AKWA9q6phkw0gnMXECmgQ5aPYEmF
5Ye/QABN+Js5G2wSGhKSJWf3AmWL/s6pP7ZrKvVUoDMUmmbA1xe35s4afsuFnB1/GsAb5S50ypbJ
pSs1i0SwKAwh3Pq9W7+L3JpGz8/MwDVqRDcWxcW6yH3BpdameAf7BCpyEy6h0z7isBbiaUNM/eUk
TFCsLJey/YyJzfPJxPQlXMwP/1KrkCJxgcE32DqiTQVqVHVBznmtkCiycv8UQVUtn/7Dp7QVtoiM
0nB/mFEzCzSl2vCSHeDawORZvr4E5rjtzN2kAoLoHkkJf489T4hjewD72rrE8CDyYDA0xJrRErOb
CjFvSkAh/oEa7RHTpiH5H0CaviEpWKs7R9MZ6yG5g86ZgWPqQwqrwRFr3kcgjt1JLlgr8XpAXJ9H
EoGbwm9NtXFdBdRDeA6V8kV7HAtCezHM/HIpieJxbG5lNeXFyj8yvPkRKsaYth2+1cdA9CnNftdT
a+2NmWuIcf99kV/zMwal5iVP4DrtvmGVnI4f+PXP2gicppxZ4OO+FvvQa/ioZY9Jp1sRcXcFW3XT
oRhPZR6m/ALeC3q1LyXMoXNXIBNFPfFOiIqPTIByyels7c65RQtLRrcQXXvu5zH9uiIj+H1St2XB
ZEWh/9oFY+QDXu/zcgc78B4kbZ3Re3bpB/7/B0Wd/ypKn9m9TLm3f9k0hQScjnpw+t+AU/sXYPZh
CR8JlHtrsh/mqpTq6NxnGDuzm/dir5ZiheO/3LDmUstjQU4qMDg360XIv10Wt3cKmIE1Veg5HtFZ
MnZXgZend9J0yDmiYCBYkF4Qfr4egOvJ/0K99w3Z+khxZojPxBCh/onw5POfYwgH83B33B4k2N3G
PbciJiuiHMKy4yEfElpwH/SQGMKx66H5ZASoNSCnEatb20fWkvrxJxnkiFEFRXL4gP+a88uuudMQ
edvaAJyRPTOEiwsKWMuQcRbP3JUH6ZHP1OK7zmpTjD4YbDSvPL78Iztqmcte7LfObOesb8v3dQxP
64dQYe4VygEMnatnB25Zdl1neUIB7D7bjkUI/xUE/reaeIHsP11Vil5a1RrJqiQ8X3iTPp7nfLnY
pfnA5U2eVS+HO5J0eg+etfodIqg66KL+FWV5qtUddg8dGqCcA8FwyGF2ORSwMB3PZvb8kXDgDLJH
zfnGr05Jabrj4+uNBxENUHoZbemhhBKC9Cr6KlFaT6tbeBVgwhCgFnBK9CK9cF3FhDB8bAZcALQZ
jiluudJ+b/jV9oEGIkZb7YfQAr151Vv7ugkpHxnz1lBzyo0jJFZjYfD2qyD6QnGnX6l8oInlemeH
zFd5axaxUE/ZCVGhVMI++IW+PQ7fMEpWtyZKUJoz+hGta4gEUsHmrej+jxj61AR0/+1+n0iyjf8a
o7d0I8AEkS+kCLoy1gwhYC4fIaJv6e6ij7/mFJrg02OtsxNs3ycSGjJj2IRRzHv43vqOjGj/mIcg
PSNf9RWEpfL4O160ILJmOkqrdToy54eMLGUcvniLlAQpXufuP+AXPaEoXcsTtn554jekKSFXe9r7
NMMVl34aQRB0W2PNz9zI/zpvVZKObDDPphwSn6qDRZs/LtrGLNGKPvWN9WYp0nLoQ4Pzj/yHfnCZ
HgSYvFQWtYpL+d+e8Ei+GC8+/Nz/+c8dlbwfEYGZ9xyZfAYyGmZuCSlJnnBZ4yyndFzRk/coHp5x
K99lwhhm3rhof3EfrDl1VeYvlAZT6oyKKY64w+xTUv449Zzfd/wYB8TGjLKmUr9A46CCU7wUTVUL
YacSaXtWqJESpz4TqWql8iim6V9rMM7qlGd84E/cQvM9xKX5hoKdE62P6782dhfsaX7pdXEE1s0E
nObZ4AkKOku3U+hKKfUfT7XZRljS1BnrefVTm7FuKnCPglHYwqIiNxzXtmgAvchBClRU6KgrtDKh
TxmyIUVk3Zav7ZciHD2mUrHmrQM57drlXINidedDpHkHRRybxRGzsJK913opJqcST1wdjHlm0pq0
Op5PQHi5xEVRB303cVwzZcMRBVzhviKo5K75KfD4zh1QLBp/KAHyHAKbNwVkD2FiXFPW88udvEvD
DlBJZWBuQVsgBLMnrhQbSvLmPXn7bSrqPOhaDwJbxNFxrlzocUifrJa0ERaWQ+hcXAiQZas4u6mi
EWrglUUXbNTDla5U3FQSaa3nYX0HuP1edUGVkXjiWyQveXnAEsNrIQA1SndJdE6pDx5ms9TePCzh
nHPgt7YEx6d/N7n6Q8NIsmm4T9tDH1AwvlgSQbaOpdaaBJPAamI01oVWWnD6pulYPAp/4dx7uPcV
LrZyIYnZWQL33W5LPpHTEgKQJd86+QFU+NDzipElq1om8fpyr+ViiowUxpHvYL9va5IrFcuzkTI7
R6kSCqM17dhfbUSikzsM5OkvUGc7DX1A3qG6lZyg0q1CA9+ep5AxgHtXfKcH1BzlIw/zjFd50Jqp
5I4eWBDGulIxT+e6pHx1bZW9n66f00YOEzdiEqc6gJuKkz5pJZD96T7aHCsKdQDcC9rWTgf8HTQZ
TFbSWncI7K0q0lt2rEkrIO8CYl7Difjh/AIdj8hkX1jOlvlE8ZWw22f9+c7sHh4Iu/BbhtVRAbkm
M3hsIKlve9I4a9HYKaLorcnrSrDYRXwESjBJd0jqmqyRUB6QoIDJxLnEfMDegs2aLXGKgeGzhDMD
bX6Nz5J/g2bXK/l7GVlnj/G03siYgcn6Hg5I1yiZSCFOSpoEIzdvBHPAM+9sRTuOg+gl9EP5O1Zj
1UjfsfpY1pNQOK5CUa2+vRnlmlb9lpZDzA94wcZr99nXMR1k9G/Ae1b89yqjhlRZ6GwVECgi4fTU
HGnF9vr4hZ4guu78D9NjsfLuBZ7tD0+M0IW1nL/pZyslyqYKTOoDYalz9RpgfIK8tV/60Hfm4pRD
6R6XnhA2HvEy1m+KZIMc0UctVV0sY0CvHwaCSM+NiP4XT5fvQNlazDiy5CFrP7Mski2rjrlfrZCd
KAxYzR5xpBViOwLjksmu6fWByKfkhKU+Qe2wQ5XP66+mNMDg9DM1xfgPph9TG+vtkTmYGlKN9eO2
eFGEm+zde8aA5R9k9GE71WmFDUhp+Kwubf7l6X2WeymTFhMNboFhMFzlsKR2s6t9i089wsMj5Pp7
TyqnVdj94oKI0b9uLVgF9Voqz6N6VDnhJ0+wl7szNojc1C2JH2zQGDUopc1TZrUZ+nasb9EUxNuy
vd9no21PJjYckqTj65oD1nRvcEGHkQ87aPoSio/530VFWZqj1tDaJBtJlADxoCOEmilBP1wO4mly
p1h7b4chHbKLQcoGM4OXXAqcrhiLxjznTIVCWsw+SeJ5+jeo54yu2GLpkKq4mvQdBrZ/NQlQlCrC
SOI5bUQngkqpo2HNMPngOip6iCWZo7pkwQs6qYuczWOZFqnsxqF9jFNr/9bLiCZRNbeqyfjt8+13
8LgYI3ZCji/VmHu1Ir7ob0uxRHbIEr7E3me1FAu6CfYvzzEtsE2b+xW9Q++MUql66Sih8S+I2BmL
rVSsPNpyggiUjfmx67L5ky8s7X2KUCPKhQAkdhdT3x8XkBDub9w1sXAb0o3HRRB3LwLs8s7w8HGU
mX5i281VTnMJSlIC2L7Rf7cw8dx7szm6VDggO9MUuQU6PRCHe8Sa1lpoh0UaKJPcpa+QIrFz6lBC
K5SvAWEQlnQ3ITlP1TidOHUZZQfZ5UOAsJac6CA6ND0eV7sLwgHnrbSVX73LBa1qXkmuvxbi7bp3
apj3vwQp036MttOKUCRUbjNvTeLfM992nJnFcJ7BbLU7r5b9yEfS4dAgFehyyUNYTpiHLs5xllyw
Sjw+0cTMW5HDz5m5j4z2oKxFUOrFrwgyoKtZQ1TPLHllgiw4S3O0HYNn5yByedY5khULUnqdRxd/
kO48wk1atf7dLO62b1IEfMlUcH9x5Eg+UFJCXu6lMTaBRfgCukNLJrWl/EZQRkxZfVfXFpNy4Fik
fhEU2Qw+gCcRJJl+u3uo7FSIyzF9JrZqHAEloxdPiIvnhih1vPdXyAxp59rWKGDN/85YkHenR9E1
TXuMN/lVQk5li4bLlujSem4Pl0NR2UKuF3cjF/bc6F114hp8pUV/Ge6xQoVRGLNBKmx0nDyK/XA+
75n0tgrgxcGO5FdyjGNGUcCtQ0S6Io9Hdyaa3MiascYf1FmJgvUaBTZ459PqxQfD4R5W19GzCWQD
2743fHcJux2x31LmYEG6rjV3PqjFkhX2sknOMvc1x1tumskiA7s6TtHdce7Fe/On+3xCwWGsWCl0
/qQsqjLCALxlwpQneigVOFgo9+9JyoY1W7UfK78eCFaVbwnSoOmlbnihRvfImO0jKUGCdSWYC3SJ
x0QykXQupvphsYlNi3CVk87rY4LKigNUObGy7sNtCv+oskfLIDFLsGrsF+dBxy0ZD5DDlX/ECwHR
6HZvQHF/NUhzGgvWWOsqiu+SIuZxPNtePvmVrN3PlpEpzWmr0wel1poXb1s6/eaIzT6/q/TdzXzp
97A7eNvsOe2NI+cyZE3QO521jMNEc1H07YX2RCo29ZeJLbuyvFyGf2/Ofjf/zzzpbZOaAu3yBynD
tKTO0bWCYZYFrVrRq4vsgy3oBinXL95BF3zGd3HIisG7WxSXn+9/WpKU8bzTKWIpXbe9TrhDho5W
jIFvr6eVN7l1S/T1YXJN19PqyTYOswr121ya0giK5I7vlzUzcvPDd4x1Kn7Z7+s46xxk6fqdUGYx
6wHRvJXZGk4n7/HaH6EN7xoCBtdnQIwzsXxU5YSifvmEyY81RPjcqu+4bWMRD/PbOzkoly2Lf83P
0WB6SPo89xVxI7nNkORgqLL8Bgd4Z/cpmjMTAtJtyFEeUZbcjpqbiEZ+01VO7MWGzLs1DtNt40Zk
LYRhnP1NmvHyTnBLNpO2RXcC3NIFKJM9kDChG2qCu7mEaiEWVvl8ua6tpzmfrmCSwsGvxG/HVe/M
2CAmsLkwSs6Yfu8Pii3qkV0eKmg09ia76KwjJ7AYzi5vQMP2WyCwBBHzCED2d3w3If2rWd2NnNIA
hqzoApNQcqFbnBYFRVUDwhWkd3Z7NT7DjwjTODAXesJjIgCQ+rEkwTLScHG055T65x70siJ+3Ays
ETFD4uBgCA5fENTHTOn3OgPZsgpXOSpCpa3EE6veToXsoTrdiKDaPDbCp5zdhb3EICUoMfAP8MfP
EMhRH799JrpNg+VFKcgC933CrHhPll9Rf6LTUQ9I3N3bl6pctWLgefalTw73bF+dA6aiArNuApBE
fdp8VeFjlZDRdVybIvgK7FwVKaE/HU4cAB5JJeO4JA4E7bvMo9gAcprwj9U4/hgiRcX8N2NC2lhn
7iLA5Qx5vL9CcKX+5nUQmFs9oTIg9ikKBYWvwrLdscp22vmWxl4WpeKMcgOndtD9J+UMEFzpih64
b0T4t4KjGzNo1t15/XMryypMw3lvS6kCaSgd2PNSJrx118So8s5kmhJ+aN8Ir5LbrB1gnUZHytM5
JhQMzVaQzUxNYIwk1eI0eRdrZuNcODlNd/VQIJEY8ZeZdlWjzusPdZZ7AZt48Sre5EuTnKPmdkbZ
cRE66xylFV1KWYPLwwKdG28Yp7/FZdykGDhyQWABtU7zA4fuHWtGqOO7ZxMEZDBPGpxcv7nWc5dV
wavEJY3l0pfI/IwgNoxU+aGoJiSnB8OodUuyFOneYILIc8rb0PnhznqcbbxBowcgWyUWE8po2hgW
wR+uArCfKLL9zG2IVQeFq8hC/Br12/16yMPq/bMlfCpSwW/MnUQ5cxTpom9T4pS6+kpE0c6t+Mpc
aKjLXk2Fa15Vg3ryCSYjkWmio2FskntUL4v8HQgQpCu1KCxF7fSo3l3ZlXWWPTp8Z9hFlsSV9PqZ
buw7DWVoTHKpoX15scFu4sPPpwKXWCyby2eUHnYai2OxGKMkB5N6cXBJ5/0iGkL1tsCDIZYSMCtA
gui6fKbjZ8+g0DmyLaOHw02xIj9VjkEeAcLFRKak0kqkfih1bxFHtBMgSAn51Pa5szHDLeNh0Uo6
BNhYI42yBV3+j2ROxGb/Pwd1XwEvyP+OMw2o2nSlAuSSJMLwM5d1ktfbR+d0sYQRGPTp8LJsNSQR
4egNSzvMTfaHKbtdFk+45rGQ6t+FIXlpCPiVT3uwvGjD37ZCiHGY6ikMapAkSHOaQKdU3kNL4a3v
fC9yl/aFlK1aERUtaqTcsoT1NdMzEqjlsAc+67WJ1snpA/UDAA0JZC3Kx+iJFWV6WG/xnXCa4Zm0
zhIm+q6T5/f/s60sun5LQ6sXKL3+SAQs8me+XwKlYQS+Hixi4STVRsPxsCVsS8Ag0DN4PLt52GTR
U3I/OOLOukSb5/hiVdNVIHHwLv892z+LMtYP0CFJy53VEhP7/q+p5PYyNp9X53vKLPsF2cEbYScp
9XMAq5MzDorUZdv+eg3zIPvvUkVah0Q/sO6zXUPhhdwq7rcB6V8wr40Yvg2BO6e8Y7ekP2fEhzrr
1Ksfue7nhw2irtFatkwdH0mNsVK1uOVg0V/3IteEB93ayLjiKAhty3MHhzreAq30XnQ6qfJqL4A5
Vwq53LnlxIk5EPCQa5dtAW1ShTgXfN+J1a9OhAESpV0h9lazvEHswcZu+tm4+GylbewyxNwk1zHB
evWVpZPZFBEieczm6MGFztt2CfpVw3+CX3S9Svj9HpYNL4EY5wvHaDylrpa1EPtsJOD0+BdrNwcZ
gRqPLS3L50Bma0GfGPwB//os/z9LCdT+oS92DTKCIH9wc+m37adm9c8oAAIxC9FFlwmh6nz5jgvj
GGNJ2pOtvKnpkl9nPPzQUe0HMq7u8bSqMSEhvBJHS8AOxxzbly50M8DJpQFMm1hcfU30r7Ts9mqN
cPRPXSHrOthVFzp+Xv7Tp8n0CD7DXH80cp1gjC5a755gWRA83BTuyB4UHeCoGKRXukY9S19r3SEw
p/d9DYXK2IMclGOxnQ8W4LPJFUPx9N8Fo0URyMJwdP9RcEm9y1Mjx/yJkqyI6xTUjHOAlmyXC1HC
qgBT3CqpHMwbC46MKopIhw5WdPuSZU3ZeC4GfT+PPQiFI10t13BtKG1Oh09nXFo9m833XtLJWMu3
/CL2hy49kmanumafyPX/V/pl3+Gc/ItzIC3BdyrRHRW3oxtx+fM5jRub0jixAN+v896HmWA+ibeE
UmJyycuI2v83a8JfZ0UUq2zs7iTi2clmNsoLNRnOyTLAJs4+4kss1OCYCI0Ev7THqXee3EjEf1Oh
DEI9E3vE1sTYMhfYuuQhhj5228Vm2kf65uTMp5bsxptTHHbCT0p8TiSGdFtS3lP+BAojqWbcCrrK
FGXPs9sZTU9fH6HaZwqKWXy57cx5SlQ+XED5zShNnIpW6NBI8ecliUqp0oOjtrJsYYT/BfQhDYHI
Ji2enLFAKNfiPXm+8mhKRMjGtBStBa7VtSLeiD1QJwNBOXSgqgG0YVvvAYLstfYMkVcgHM8EYarL
XGm4uDvfIOvg71dwoB7XvjeTNKyOiNa+SJkr6lPYO3HvsRol1mWcCQ87to4zK6RgMbo/5B9VJPSv
sAdtPwAwQljo59ChAJf3T8COJzYVqGxhacpwszxqKYRTAVHBxQRiNekzCA6D/N2D7eEJdp5qYPyH
gnm76oVr+3kfkvWLnoKQJL6Wfq6itSlMcphbrbC64BHo95sSJk2mepCikPqDML7NFPHaj05ncQvg
+aPCBNF2STM+GyZWVHyEfYUg43lpmhlqRvhl0vvyFT0wUNi/8l/slrFkQKQjHE1NGwD3SF7mzTPG
h+O0lPhwnFXQrQ9PXGQZ9NgG/2SPzI9UiNzlEnUW4WqQmWmHSttUBMgdl/vHiIbJSfJ8SJODXW8M
ckwyRxOn9AA6/O/YPpQXV306iblpUJ9XNXh+ygh1LOzvpduGSVC99AfXqotGbgXAIXYYXcpCvEB0
gNnWH9quOZ49suDqciLV2BZ6W0/FQ0KIlLeE1Y4gP7bOqWbtrSafd+WohKZNlREDgeuXudVYPqjn
7s0CmbCbi+Kw/lAMVdfpUlXkhzADco7KAPchDqKh+h0pO2zlQGiJ9IPfYqp11URIak6+vgUazLxP
H9sMtRPTnKRPFg494/LHOVuS94cwrTP4xyE9gJNHLUCIjxxm+ConS/XnuHh70WNxhKe08IqkLhPA
8faey52lX6VziHI8BxptC3xYdBO3EGQTjJI1PWMcejDsTgN3zhqd5jdMgGevm+8wETize2+u8dR8
SDSRvhwRzdFbzuzByMpXYNPfr2xOgkniAw8qnkX6C57a+/jl7SzV6ptGIMQ21Ne6IrIX2qpPhouQ
uEzMF/VxhQ+QYNfaJtaaH2a61/6Nuy7nzA5Nv2gwFvyIdx15ope1SFTiT983BF+FJILy4SwanHAw
DYUejEZHzte21ZrQABzKCBAyfbh4b9+rQkHETtRCz9L+QrdkhQuMs+oBgAwSJ/1bliTnshpqOxrF
3hLVHGVP/M6d9NVAXOIHqss0A1NrsGThh9vDuUFYIc/gNFKBxKWxHIBXLo2RzGunaF1vry6tWBEt
iaTTTgNtQJTiS7uux15PUkOo9VvBfN4Miq9NK6Q2LII9KwFkpm2rqfxNJjao9rY/9DEQDrYmsEdJ
B84RAvInTU5NSij5P5AqetTpgA7JdM7i9qsIxN5hGUldbOtgEHog/2x8VIzm9fk77+34jv3kJ94i
ulJcyZ1XNgIHZzJcpXKD6OOB22uZapo6oOh/Y/BwccPBGScPLe4ShS/k2A6DBwBctMozuye4Wf1I
en+fMJMMIBzY1fL/NbfJRTxJxpaNE6kzqxnFQkf7GmeoGmZdWMSCvSFYhBk3Lk4j1oi+fFLO+hrP
Jv7RFD+h0GrRhZsl4tyR2NP9dLsElC/9WUlfUv3MpSWBOFXu/YInoAHLE53MpGVj28nV4wUEYFMZ
zzX3mDRdFEH3sYllc/tQtOu4TImIcY8JbFydqSpUajMaFkTcj9MrnKDgZMdBkVBhOTSA2Rf26gvJ
rwQ1tFwZ3JZN5fbSbu/HMSrvXQEURqTXtgQC+03izZF147VR7DIeZcu829Fla61CYm4CzXi2W0S0
rwsXL+aak3JOvneM2O3z4jQM+gkCPd2KlcioPr+RgNC4O6JEgyYoSt1UZC9/nmmSGhEMHfSf1hus
uHJLqcPaO/+GXpDrWJjdAq867qVo8jPDsuhR0hQG4iN/zkTq66uSMm8dtoAJyED82hkF374d076f
imd78TlWPd5oDgHXi6FVIwD0lfZ884yQbp9IEaWxj5doUe6B9cIAKfubfuVq+VojAJOxrtx/vHxJ
RdCeQYX0nrlW5ISSVJc1ifDsojNhZplolnx4j/bzIZ7LPBJeCZJlf/kE3VvZwGE/DFy6Q0rfvox3
/45ZyyolOX3nEo1/QDHar/sKHIGQn2v3xUxqovLzSdMjE0IXVPTuiyVRwP/TaWtChfF+oEaJum4n
2Dhz+K+m49q/eOzyUj2AFeT6mzyJdwsT0YzYZXc1KkfZhgM58Lcsm1hR9sRBgiaoB4rwFwS0Dkpc
+uGOGaSmiINYiHj2IYFMDmCf5WlKWAouiZGfx6LzedrrWZhu/L4wiWuutIXMM3RF+uW/Nz0E5o7F
AFfgxBEkwbhvlgEsO5oztVHR6zn9Y9HsIrAn68qP+CKYgDHOeygGar4o7eQcY3OFDnoZyv6f0dDZ
ZXnUdUezs3x1yM6G2CILPIfcXw85UfcdlF7DFKDj4JkNT/wqJi2txY/LtUGLQTzBDfbbdeSOU/wQ
edQwP7meBq40Kzwf69D9Hm6ImQjv8IUld0ndq9pNxzGHZ7LDgpGS2OnkDlolJ4e0f0ZLsncounac
yaSWjJW5huaj58uhxfh9b57AAFo4bM04cKs0AWpWDzzwm5ha7zuq0pBWOu/jbccrs1nxF2sskDoi
tEhYotbTX2rejk0AxEX3WLwbuwkw5v8gE5dRSdTklHY9PfsbXYcdAWa2vTB3aVvwYjeO95Gz/in8
xyu9VhJvWUnmm6l44+Y49iXsVVz0Cq6GMCZ1qdFIeUl1RK/Oyrfd08rFxMlOYXrgSzs/tLFfti4z
a+Drbi7UoS9fJ7KoHXnslqmgJsl4cCK/Vl6XEl8jRNThW9BbQ8m1a/Db2mZZA3S23NuHZEZaVw6f
BnddLZO68UUe79gj6bM9uWQGmkZvymFq6i27OYemqQ6G3S3qtDrpYoSZXDUKh2ftvDJUu1gsxMQW
cYbXE7OdLGwzEcVlnVfHrqY8LRZZA+F6iMGw2mHdBtwj4QdAGsO/6Z8uIo/Fg/HHc89v8uu86J1h
CWNGaQ/+mJ3+/AezqHXVhBFPymkQSWczi73CpgbjYi6tfKNlC42e2w30J9jPdhRLTxx0S2B/fsT+
3wv0fs19qaFBJm0FuebWRdkkinUGQSqo4yMkwWsRgWB78/rf3H+JWFTyekgYtBCq2j8VPrPRHcMd
JRLoJU9IPoWFTHujP0CQAb/K6V4/WMjHVxAaQkumtkNiOPqajDyxxRl0WbFaN4XWo4U00Qo3YQPW
Y2Yv/OviZMy2h28AROC5lce4dioq+Q6u4DACLQLuwsAEND6aWnQVF06TEltnsLA/kHOo0dzP3/bE
NjF1ypCGLVuzZdiDPySIuip9tyHjdsAvXVqEV8WOL9VlXoltWBEDPYtyfVfcBkcKBgC3PIV4ztLR
0trVhQNzcDGO8cx7X6Qz2rYIBTVxKnVMV6bLQeXO61y2iMoen/PTqK5zwmfZJ0dc64p04mykvS5W
aGgOQhfP/CdEy0uCNiuu3nS9TefGlL4DaN4oj/lrCPhw6xiDq9MI+DRbbKDQuPZ2DkQaU4OAVbXJ
NSBWOeiM6n3knaTBNxYMir3EX1xG3qkUeO4PnbwIe4tEMlnod/1ZOsp7LYYq4vbe9N1Dqu+o+a8D
mxr3b1uClDZNFiX3ylWkqayP5oH3zKhqHjqI5QPKzTyz28i+Ta8c0DS+Kap19wnOqhYOo89XqK/l
bf4hcA/92/qLHnFO7o30DsETktdDVISbb45JB1PDf+6V2h7gnCS8vqVp9r1bQnnrsS8egdZyaloh
kHaWCeLNLe9xodcgsYu9fPY58w/8Lnrvl0K18AH2YSu04X+s8J1ADp8y1HUxMC8d3Wso1tpBqQ8p
YcoUYCD7YkvjpRkbRq5+jaXYFskN7/lsmgzJ4Xyn0UGInrb9MXMbNeROlU/WPJumMD3wBdPK1hpA
xBrKOwSPZqWR8tcoK/c0Eg1S/jXZfAZENmgWhuSPCis8HsY+D11UTLonVeDjySw3rt6+DnKQX6Mo
LiwSJ9ujsaTnJ3SjxQbab/qacZNR2ooyI0aEiFtc5H5XHzo8oiXqUSG6bG4P5xVsQTQ3p6c08J8P
SmFZHZ2rcZnZjhow+7C/3w4aVEYioHFqZSYzswktIjgM8cUWwxDfLppIAzXaH5jfj+FOTxXu+Igs
cpb118chy1E2PRUeHnsSji1xGJsgeOYLu2XPR0wViMznXMA8WY4hw8uehnRHeijObYPLqUye15V7
JOKWfWqp/aJgMV1hQyA4xGo0MvZRBOdln8q2qrnXTHeF02ua4bkaimlx1OwhVsNySX4JQUg+21K6
dAXtd6kkDkeVFYe2aygSApG2PPvUPTIkcg+9pw8JFu3RsBYl4MnmbAyvf6qQ14XjMTZa63nYyWq8
OA8Ymf5/cagSTMjAAhn3sdJAF6lziXxotetmNOx/DmlcD33Udt7N4OpBZfW10hbRwBOykx1RarJ5
X8AaDMZdfvCtHJv5g+bAK9IkQFb1WeApp4YaDfu6rSgjXKLR3k8WSuVaL1AsZpnvVfKdPcQ35Ajx
52+o1Swsm2s2rf+Fb0zYs7vPwEbV7XQi/rh3Vx9sWL9n52ogNv54pzQEkdI8gBIirFHVeL01SOir
AA5c6Swy0sGIn7hsAkHgOFyst0gGoG8rCkF1xJwLl6SXDmPVj1kQPVMYvUiSlu3Pa3raKpMBWwc2
SYTwi/mwMMRCfgENls+OEB0Or9udmCyCZ4FyWdLpo5YETkL/Ox1gVKkoL3zLPL4utbhLs6d+vpOv
7OhkUvTWW6R67T+IshgjXz2yY1Sl5/k69AT8Kh0oyo3zoRVHR98N6x/3GyFKAsgn/t5CVsIdaYJk
pRB/ZnffAvKRcnj9cPiMDeoxId8oJBDb17/v1N+O4WBDsCO+1jMclV4X6L+txu6hPFmtIbPD1yuv
DaH2gxcKuRTfMhcXLZwOYmxDHLP27XJKCrhD68lRnb4MMHgnMyeuU/gggpYMr8Be2tHyT0HYIH9/
8xKGGafGa4BerIGxsbgpJL9U5tJR0wsY1fTdlvJ+wSMYhUdZeVpVQM7PUJV/2CTrbtCEmQv+LWZ1
Ionp96Y5opin2VKANwONaQma9gLkYhKNQvA8oLmiqRps+Wi5NivaDg9/N2DW1K2KtZ1U8T3mi6Oo
Oee5nCuK8NmaQ4hflD8WtRjxS1Th1jydULRvVaiEnSpfMfez3acpjaqU858KU0z1zBVsOOSzDevI
j2YKC+ZYAC//Aa+TnuZfAQEAA0DCrSS/S0khXljKZrnBrpw2i+EfRHcBmo+UnaPGj1ljlY74u2d4
weddoSlWNKaLuzzzCOyGzigRo/YSTPpvPBaZr2ZS4twbjqrXqz1UVhR9tc8LPKgzky+KQBCbDp/N
zCYdsxKszF+eeRfznqBIx0IZ/Z92a1oCz7+JcrSmT/zujqiEbJxebzA3yJ/yZpE+7HYH/7AqaOMQ
Sv/UiAdt2Kza8EkYFF2QxxQaBYjb8fcSK9HlifLLin3wMoI5TEnTVfYIKMFWcflR7kIpEy5k+8LT
a0HfI/MULDle5SGqyvKiGTjNGDuFHxH6wQVP4DUIYXtRFaMFywgP40B2VXrzJoMgMeqH4Aa7rT+K
UD0OHluK8e6I25HqoUe0YzGNc9nrM4K/p0eVakRisZ2DVY0cOuQKTA/BVvIzTBQJ5cNY7h5E5KsR
ocagT8kXPFkjv107K+nxKGJWg03aKjCL9//b+RZ+mWX7Cs02RbgkGnORr+LV5p4K0AH8WN8YpUmf
ygA+Go4om5Io2oibLaF7DsU8Hd/Cy0EirtqUVfzIK25L2yn47p0z2ehV5DENwNb02aHv9igquEDe
Ca3XpKZXlk1IfYltdO0eqnYMTCAAjAg92v5gseECjnGAMovqfn2UeEPGcEDabZXM5kixAfZVQn7n
2Vd7m0uY4OkwTYndtM3/x26Eq9Or2zLDY9aAXttIvfQurp/3E5JSIVsACz7sidJjcgntgvhktZpy
zoQPXRoFGW639HHwRxtubLqLrVYNSaWM7aSgMLEAnxlveueFTcV8pRBtebxzRb2ATLLItMJ4PjP6
Cuje1VLtBVXlLyNJ/k5N3IcIdaXF1eavOQ/suFZcoop5EMyThGoE0HEeZO7JPUf1+te6kfoASj7S
/6R/PlZ1Sh+RNWqcQ8ggrrLJLGkTAY/MJF5L3xMTLym5CcBvA5FBBoOPMM7HGTHxemhTOQAC/KqB
CeRqeOYigmq4JJG7Xi4GYrY5JZ94XB391g5lkP1lGs/dS83nvjS0SRVyH7EzyEtpFm/kmzRfZ6Qt
pwIoyq5LNo0n9JARGltfZV6xGeqduiGEWwN7oR8RVHudii1Llh6CS/38kRwVsnMzYdOk4iZJyIpc
bLTe5j0OJ9yYzo7BCcgyEH54uYETXXNS4cP6oEH3gMlp2aTRc8VQev2JQ8CH6zc68gcoSVOe7xrO
e93/x5JQw3CH2FF71CKEIt5P88y9vbpQX2nXLoTlLusIfxpJaG+HAvboxPJjidOqF+94WcCubl/k
DLmlO/W6bbq6CTumLAbxEFvIrtOzHBkYhGhTrl3aFU379EEKhVa1Ls4IF+rLhUwS389Tb2URWlPo
qu3W4UdbxefxO/I1ER4oce7NtqCxOiXJs7howeDc1uNGd7Spye1X1LNdo8kHmRd5wf9g/P3HQIKi
U1Cp4CIpH2OzYX6kqqOmQEmSX177P+CMVSnG83iuqwA1Du+l5Db3Efgjf5NCdkGsjv6vo3dXmdyz
u2E4Hyx1ayaMV323D/3TWEBzSz07ZF8jU3sgvHeKZnuAp1Q+Y0uUK1QmWVq8Puvag/aA21Td6LM5
qAwxNiosGX75lyhD6vn2c+2QmXus9oQiQsKq4W/TtHvkbLIjYKkjijai2Poz0xaxle6CPyz9T7i9
kxAM9VdKIbrUozPllcY3HsfVWxu7RuKC7JCHgw0eXtIkYicoy2z69j+PrUgluiYVfxfbVo2l4VSm
KtIn//h95/B3yK4QRdptc4R6X1imPCqG0osx/JuluO+0Zj4aZxajhJw1FFu8PWlEotcAPH3RnRjh
/WVT0RFzrepLkwvl7JXnwjt4KWuVQAvvmrAjrxiNaD/FcXXGpBX+p5mn6KwW0O+/kAJf2ApOchee
7YyCyysY9f3gUi4ajiES8T6cBqZseBBEVFDTQ9SIzEbgMH8hIp9RaSrdthGamvLndylhmxBuGnTE
GZmPEqBbE76w4YxOQrtt38cZ/QxeZ1yrFCZ1wmP3NMzn/YtJXnD3jElNJZ67IrQInoxGd05sZKr/
e7XMM4ndTpEMhx5TtvNCyrujnBKBy3tlNwnNpKFL6mQEWywWNJiOPbAW+p3pRPGGVMn61escyoCj
skZsPpzLLXqxuSc71ESuqB8HLEiozhuHO425vb3gvEsLj7rsSNiLl1VGkwPdLURpSf+ln6BeTdGN
CHszCGfviBQpXnIYCA2uImPJHqHPLWMJ5bKqwWelPksREkD5BN7VCM8fEjhBQS9fDz1SPaBxSkvn
JgEpw3GUy0Tudee0DdNU6m7d80x268Ams9z9MamRudCutwaco+qSDpmuabncLZmsk9SK/RlMuGv8
LP7OoieTT9EYaYJkB4gXaeCmdWPLmgcHweWIH3DffIOloVJXjWc5E3mV1hHAgdgyVxQRQ4y6paiR
I73kfTK8VqqCoZNUtPnfx3YHS6hxAg3L4zwleNOVTf/DVvcDg8x25ZeE+xCvkOLb+hQStKb3KCR8
9trI08LcbjedVoM1o7Hu1afrfXsgladZV2EXu1O1hFPOYAuMxi7GwlXirkNHFcw13uDSJZTcT0u5
Kuo0c7pTGr/E2/4xOEyqJIcJD0kozKC4Vh/ep9IOAQW6TM2hnw8/TVSNAiMJBXrulKbZrbyu004/
3B2tFqg0FClL1k4J3qN5LtIKuwQUjKZeR4bHHipFPwBRon2cfBy2cztORCOQZGE2hVhr/jHWkTu8
/k6hjryl0KwuFg4setkTBaB86kGR1nzhDqu0UD+cHBEsCvwkuRt8WgcpU8WHn1Szw2INcqlq+IfQ
Uicm8VION/4m4+KxsknKll1f9Ae+1HCRMaYhxCVztNL1+9VS6QA6R1Cw65S4F6hAHPXUWbMcBfSW
SfCO4eFV5lfVrIamjMBxKJJOPdLdqvuq+tLcaQJb5wIjUiLgnGCoCfne8BTrdhrkKBV3gfu+7fww
GSv0uhgZP4rv/ORiEjv5vxbBu3mBGpRgk02P654A2OJ/l8yINZoDYcwdc7pGZiD2eQmqAlNQh0q2
fIbTlxOMEnApZeaL+PJWKY8B3d9rdmEzWctkMGq7P6D1OmdEK5ZX2S8w6mvQiN9UcZcSeExf1Jbn
iwIuoKMHnAmCqaFUrORaVcj6G1m/uV4BykSI4Fw56yRGkX2h8NCRQveK4PVC6iTe2Q00rfqDLYKl
6xXNonsCaOah5J1XLniE2uLJtwNppLknnvvDaLzj8SelrPSgm/SNpwNfjaGjp5aRekfrkURBuXt9
2lCs/wfXCNNm/LovQg==
`protect end_protected
