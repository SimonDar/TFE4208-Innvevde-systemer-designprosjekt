-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yDNzDB71Oyb1O6SqtS0HD4TiVyTFuZjqQfPlCuqxfMpuj2ViyVicHSbWA+ObxbOh5kngwJSN/And
9WTuyZ1GOYb7O0B8cZA632qbx9lizxdGXO5h0T6MF34xW7OaVJQYRDe4aA+8gKTVO/9Q437vz8Ff
3O0UAK93c4u/y98I8s/UJ09Xn0bc8UtC9IKB1VUxEMV41/AjXuv0VS/u4a+pPoY2+2R+yGSmAOjX
Bvy/lY1EUTNbUVxzmAMxlHj5eOHycs0QeRmmaqR8CI7/i4EdZoIo3K7WdFe3Ra6+fIjFcnH1MFdt
Ku9p/HkNy0pTwurb3cPDJ33vJRqp5xqna+F/jA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
vKaEODP10BvNXvGQFDyw05uw1ya1pclq/+rB0lNuXles+LRKIW0XUsZuqYcHqXkbikZ8HU+O/L2S
sfFZn6ldn3fMmSGRrdaF5VIZpJgUWM7P+B9t431wRQ8Kz+hKHFN1KK7UnchbUXrDlUEG3JF9fWaZ
8GAbXMGviWUhz3xbp5WII3byD/+PcJ+a6Z3EQzUDhjf19fwV3dVmhV0P0gYOhLbGWWzBnw1QMuMB
ySSSX4DZMx57lHxpIpBWcdVaBGohh2ntIKP0LXvqcg549x+b/JuxGhUBrN/0Xg48NT43qX99iBmy
ZAIbx4LD50mYJwE110wVv+5Hui5p0nnkD+ZJE/SVJwFjXI4FqTXfFqJY/486Qp93QzaaDRu2vssp
gtW77pqqEsXmFyU6QvQiNxuYZVR50aprsnJEWTNWqf1DQbvHfDNJ9heUo+PsBx1JPTQA+97PVi69
r6lkSj0iV/rO5Z3xbJpz7xRbE+JiuvQif8VRPkJMfu208x8vL/D0aPuLCxt80Ekhv/BcofLAoPpN
1gpIBz+oInoIE1g11TFo521rCtOfJVsbVJ01mOTMtIVtN2oR2o/BpZnpRGzDjgDBotcPhjAZcKz6
ttxZKK5uJPAFzQ0fIka76xwrcO+m+ayAsUQDmM2V9qXU225x1EZ++VAlqCUl+QC+oKT52o0EBmmD
SPYU6pTzRx+IZHF+AoRSFzj4JQsDK9iIPl6yqnmQeldK2zav7O8sq5Bc7EnZTM19pVwJsW+KDEWc
/gjKP5C7TagkRXegjuRZxgT/j1QGLy+8EHFbP6LOoCitwJ6GZXsmUs1V2moB8m2L3eVIhdG+rH1w
fitWofBOEtWK6VPPM+7Cvcc5KbUxpFfW4uQtt0/S3AypI8UpIZbel/w9oQqAKx7hOTFD70vev8ai
XlhhXQOR4cbAmz3lC+maqkQVwqAdipkn5A7y9oEerlTeClpE87Xvf7C6w9Dtfvl8nq+xXbyqclpZ
nbjmPZ9fS0IW1S+rZO+rqSMQDavTR+FlAObHJLAI0NCTNEq1wBwZkr9BBejwzm88QBTHwgSCy+Lq
kyH7rvOz63wY/JFCatp780DgFs/aI02UmeDgV66EOHS55VXfaXnijDbtAZj4EAm4OURcEyc3tiSZ
hsnz+PbtWyrSss3NlXMs1FhbBVGs3EusgQMz6QHA7LHA6AWukQZ60k42Iq0t9Oncc1ZpJ8IoFqYa
7lPu7cBiCq/Rc0qTWC/BBNi+PSGvVFix59+iYtxHoarHy1Ka32Dtl8d5xcz6BlbkSEvgb9NVcu6J
0M2S//VLU+DHxgnLFujkvFCUmzSytbXB9gbnyvGuTHIWt3ZRq+dWa/zEoanOsVAAYfzyM3sylB1O
U7sKegt/Zruyknhz9ZEmnn3fQmTTj5zb7hUkFoMqUqlut7imk8ojzRt5cweT7ZH/Pze7tTI2CPKK
Xd2SuECmeby6ThpM7I1wcx7qANORsbVoXUr1y1ODyC2NvqS3U8XmtDF/V8SbxY85PG8+3ovMYlW+
lneEfLj0xbNLWW+tW22Wd1LLTLjH12Shs120RlK4k3KkzGD58abCsvzdMsQ2a5KGncvaoeu/Eaph
qW0dt3WC3WR+g+0j0MOxZWVu1pRz0L15F8wG92AKDIveutqI4LECi6MFShU9G3327eVo73CfZUGK
Va41i//UwZMsDO+m8NRlpbhknTY8I9CO1P9fPzxvIp56VsTzuz7/0Q50YvoW1Tfn18EWTB5xt36F
3unG70YqYkwQWTCWrUWe3/UwS3VNx7g3h/69mi8c3vA4US+DKdi0NI9EoLrQWiu6KkgfeiHrK6kI
zDk9lMG42gB1jeTnoUxRtwOGnUZ4ui4BL3d8cWhYzPbM+V4mgADA6VT5PIgZJpIjZSRPKoCMU1g+
ttTTUpAJBJzfwtmfyxBildGl+/gylZ1E0ouZE7nYEPicW7PrNlfFah1UgEpV+6Ce3KDfCPJ6AjOE
8M0Jw8H0Aj0z5enIj2FYD40UYFMDLp9cthGaeg5TAIF5wAdZVP8/FJGWexgWrZpptMgV3gfWByD8
2420CPDjBF3+F1te3UCqalb6xWnCfNMR0Gd35RFyu7ObcG0unX/aot8ruK2fRVY++qNP5aI619Mt
ddSEK4+tPr/3LQd8jbflYefuN/YHvtorgH8gsRN6DQCFUv97naRkFjmG8vh/Cz9JDfgNnbC2bRJn
dYNy3TySKpFCvCo5hyW7W8RH/OWWwrbv8FYSYjl9HzLpTq46wkJi2vIh06Px2Ktcy3QkVZmMZ/PU
tvlc1dKSiYZW8czEe3yLaM2ka41VvcbSADn3aNvMIAVDSH4AY3dqgYkDgxpK6I5GIdE2FEpsHEFA
EqUtdRfUrXbqfwLEX6w+GPnGKZujy/ZkjYHMY/nYD9FhFYRAQD+wbN13wOmfykKpf3j+SNkz/eIZ
pd0n0F0hHLRUDUcvEEOKkrZfETuAmtMhYgL3XHTHsfDNxCb44GP3tW9NMfq2VmY9xJvRNgoSaoCV
A9XMgMcMgipk4uDsFYcjB3Q/c+UBmA81/xHwyCvhyOM9P4qDXZswnA5ZkFKKJmrizzBkF6S3IRhO
dcwbBItUlI2ceeKnZEDKLmDP7rXect8vKKdVbljJzGXqI6LViCRe0lFnsY2p7ne+PhCryFop2rZ1
esizOMkyqloF6Bcz0wLv7QklzvLK/roTzZMz02aZPq3qUkle30atf7hMaQzyov7gtVOwMILbaYhD
UUFxdfsAUv26nbgcNtXNgYWV7V/2UOwuZy+RUdP/iG+K8GubjITXBxygOEmZ4il2sxl2wNZwe8MN
t0VwlPACfsQj/Cm8LnJekfxSSra68RcNhl8byxBwe7Mi0Lr3tWWovuqw6nO9B05bC/BQqpQpyqQI
jeR57S0RpIemtMbFzDrM23Li7Nlit9Nu9hLJ8sQR1c7xlm4o7upflPgjAsmXRo+1X62iOo1NW5SE
Y+4V1mA4lpwVMky4BAjkuWFCnmoArcS0RGEBsXqlyP0xpCdPf6AuLoWIDAP5sfQgjFjhH50jxAPc
tm5VIfBVekCRD+z71wgzMCorjUtzcPurt011iTYIUyDda11HSRujpinasU0Cu2jIPUpv2evO7Ypk
bQbWnYQGGOltTfRrrJ+FOy95R4SUVfU0WqYt5xfKk1s62xpnRCXwlW0h4iu48Au805qNywaHYN32
c/N3imO7cDFRWEP7GVA1tMOlVMGiV/FpjL9oqcBUYRBwRldqBbenNL0O2l7UT1K++knL7+/6WlAq
QqMLxEsG6Wn+Q81wFnJhc3k5+9xfKUr7s76o6nl7+6ZVkQdWapVHzCC9GYOzRkiXyhVQ5Ys7S9mO
/Go7L6P7BEzfmSNjmFUQaw8l6eq0jLUwR822GB2eEaSWmOV9QBHu0VpFJwvG/1D2h7SdQjuR+1WZ
x641qVoAFB4gQwuQsBJSHgzTo/HqN6NZS51YUQjjEWom2666KE94NoDGQFTQJxMHT3vw84pB1MTp
FjhuzFurpPG3gYeZGAOC8BwDzJRxH4JxhcTcA9AeV7ZEb29xt95rCbCX8kA7ycxfQmazH502/TG4
xfitfujYGXctoJdGCZTNaeHPWYUOUCgrhk5OzZfY8ScVNgILpw7HDYeer4j7EFLe+wUshI7BEjFD
HJBChqia4+qxq2oTkmt2WkpEyIx3qK1Has2W1q1Si4P5oT+Bntkcj/XSBogHYwz0E+7nX96ni9gy
kx2mK2k+shBgdcX9Ov5QPg6TaaMElLKYIv/TGrY48KEsK4zpR516UDQ5s39v7BqTotSWUfb2qbD3
CzCgH6OtnN4IsR1RmMEmY6/cZ5HNvHAgu0VCcNTeMZLMAV6JFcf3QI1wfjBfoX50sFC/U6YHXMx2
FnQYLKHxWsoKr8S2rO9knuy07xSltMA+2YJN0b/wBi692zevekuNqWcrusncG4bQgb5ApWk9ZHpu
VE/3rT3mNEbkb1aiIMHA+JF7u+gNPMQY6DWQKdDBu2Oq9kI1y25Yx10dqeWCde9iLZBvjbkwjxDa
+hoV/Q9fN4qbmcErJdjYSrfg4K2qE96+kWXOL/4GcMQNuGsxmWXHgJyadh/V1PjyiPpmGB/m7OGN
lrVz3hyrajlcyzooMFe1uOoDMm1Fl827/zAZ7lJnBUv+9vFTQ8LZ4Dey9TsjbJdADsaah+ll7aO9
53dZ7/TGCrwhPF0OEZ3wje8xJnJ8xtQVZsOCQZjdpLRBh6iRpo2N4JFxu5FL3iEt/fOlQO5wkwja
Rb7bRsDHEfIVvb5OtJrG6yH1m9XvDZ5KAhKLyJTXxrGh2DIjojCWDDaUOtLLbRBdbZiJEZcwoOzS
s8BMKNn6+ic8o55IILk/VR8QvJyYDwtjz2tsrEtAnXYTdRFmQIcgaafM4LPn1qX9W4DfffLzi87Z
qT0H2EvBIsVAVbK04RKpyTB1XpAZBMZ65/Ol2sTm927OOhN2MQthNEFXJXX1T/xfe2S/xbyE21Zh
LF17muMkRhLja8fWlJcx0FoxLbXD0ducTon22r4/CAuYywsnoGg4mteuEY9XXa7f6dFhqGyf/D/Q
Kg+JSATSM+4djPF4E0pi/2mbKqm/lLH+p93sIeoVWFvGRTyTPVRFMmBDf27/ktbW7UlMWo1+U1RZ
ffbReBYQcn1xLQ+lWUPrDXWE+OM9OhnqT/gAMOACoptJ/6odWoKaRUmaVSfdXOhFnWmj0xZ87gT+
RccAa5Cz6F/IKuI5owvFiIG/VvqqlbKH/uxK5nK9wp9Z5ZAOuRSm3BtjwG1Nx/XRILWaUX0AiSET
nPj8ebLXPSavmPNfQ3vTsMQo5JG6CKlNQDQsAemriXgd//uD9CiHEcDmdmxBjtc/oBvsyceuf8C+
1T9L6ExfPQU8S5lO80I9aTu+CljXbXU9lsz8WVD7QcfN8Q73/mF3TGPFzoIA6Gq17woY1zWxtWUU
ZcBKwdxTUc4NwP0UjSXQjAhnKE9EjAfNNXmthNBDugdFrvkRiIY4Qm9gndCiirezRSSCQOweWifJ
cjOEZ/7BOthHq/j5ciN7+7qllcrrl8B9CCc2MPfa3QY4BeXEdwNeqrFywCU1Mode7xP6pIc8Xa9K
+SIO3cWEjaLshZ/oLWnjWt7/y+2OShAC9CDspRMqEXEnkhUKCx9zz1uQ8ivO5++/mcilr7LZocee
3UEaHWe1SuYXakw6hfH6+FnnKe0KdnYIIkPP8LntheBaLOXfj+PkqlzQKFGiNZQVA7m1fklW1Xob
tcNn9vWt+m0fsrcUqGmto7aGgd4WqeJAGEjPku5k7VMY4UXG/k1KXWrCtEAscmvPe/WHqLNQ+hjq
5bTErLCL5JG9RMdBZGfO+JEiSC3TLluvrKOOWxssLTAS3FY3XnuVJbKILowOj/fT0/mI8xe90GXd
4rxBcfZrCUGhKlL3H92OBfNxypROCWz+hee1Pq++EAu/rs2BqqUzzV6TzHfBIom45A7tNosUFpZY
c1qFzqvW7LGJoRkUYbSszIxyBxPYBInrkl1+v294XA29tfY8r4oxiCp+RKVRLeOROnWD2NLwdJ7v
GFd3nfe2zfGCjqGxxnSv9bXegEeSwfLabISkzIrjxD4fSygkG2xZQwCDKT8OsUYI2wofCSjR6Aaq
Vi0s69/XZO9yeLtoZb/Ltzdmz0StQZNCfzrFUOOKJ88RKdhDt4QOdXaWBKl4WDhTaarjjzUgHp6n
v9sdxSO1I4HQJVeuJ6E4fDQpjKyxlHEAitWuwm0ROS4oDff7QT6Syfx1MfLWCm7vR2Uh09856ZDp
dOCZX3z/sSbetVnEJAclghyILgq2sGq+ovoUVzyyjnyBFgTIrDpW5R8AxuINgRQj+JF6UngKBDcI
TXjZRsdK5zvkdTEd6oaw8MNDVZU0BFYDMDnU+gQUTfyVCbTX2EnX9wbpd91FdE7AgNSmwuhRsWJT
jC8dw47DpQNix6QcY1Gd9ba8gh59aUz+LyPKSRTAHD6RPiXxytd1duNKphPxRI6z0xR1p7NekWLh
/+nmbb8QzpO4b1706d5YxSVdBnGr4Pg8qusekGQpmQV/Ub3MQoCpFeGCuuMaDXnqxcsEKs7sV5lb
3osOBuGYeLuywdYCPUPu1JGSiZYCom1Y0KSQJUw4qkUd6L0zs5zggWxwcVQvJTFlcyBfN268FXFL
2/6jcdjJ5px/J06mERzAWCubm1d16ntJFRXadEq7r//oEue590H3gMwaQk1ivuxtXksRV6dS6/24
DdTXgk4QJ0v0sSHh30z6AoqYTGdHk6QSvhdQfLd6JGucTm/baPc1uURlzE0NkqEY5w9gc+i2LwyM
2R4Vv2Y0Km2+H8yYNgj+CVuzibSsLZDJDD3aCW77S9wlKnNCvqYgTv3J5egFE/6HkErk3ltE6xxz
meAxsWf81+Ssz3oiD+cccaOF2cPH4TuFQT/PrmdwrBiaC37INXySkeCw2DlLAU/bQZEVUjrpK/W/
nCkbI1hERQQvvkY/QWJSo/k1h2+CJt5OvjMc/2LzS1ewVYB+mPftO9KkUstvdvZUwKRUgAFFluYi
6z8gyDsy/Juy56fnfDeuFDx6UiXX8HKD2Jmpb7M3uNVL78CCDk5XSurm2huoyx4R1lqajLd22TcR
Ykh7u37ftvhahK9I04ZGsrJx557JRJoPuF5t8OC1WX+aiwk3S/IpzWGuZcG+DzOswv+BfLG2Mhzr
nC8iT1k+9as4n86VzCEynr6qNvKh4bUj0I7fnajcDUJsNHEyOxGly3gU10h1h2s1WSAwr4GNyPs8
WHIfvWhiwdS42vs8GqSN5b5Hp+i6oZXsCq/05sCR8ImFhtJsuf3MoM1xRKkP+/iXAQpe+j4VVzbk
UqI6SaDvc98HCnuDQWDq0cGdhgt4BpgPg+48wNDCIR/5lQN19DyNHveO5HSvudVzEi5dy33valWW
eYceTPWguseoGABq5GqruGjjMAiHR37lQlZu479phKNP4QJFotXXMP0vt8LdQDu6XeiHvBA2WuBH
h/NVD0xyFPDEH4zZAT5C1xtq4/42eTwsqes0Bv20/2fo5OtXXRj+p+Pu6YkAsv16OYDf6l2g9OEV
4S7AvCRLktzrhheGllh2T2QLqUQn2h5C6fLiIZJk6lZtomJHF5FPXlJWusEWKGiQzfRJqK1uJCjr
HVQGnyKyENys4qAxrXmWYrIjpTWYfrAtYS0Kxc3XH5Uh2ptSL71ZYmGZh4XGoXpf/0GrbS047cEC
DlZWNPUllvrms5bx0SvBNXmGRRQ7z3+heUvyNFY+/0I96R7KM49+Ohyw9duaNdv1VU9kG7ERFTbw
Tn4tSe0wcAUIpDIuq6N4OvYtm3C48oYivx/JNnpoCoMk/V9iI/qm8GyNxGNh6M+kjn9a+HQQFbUx
zByP6FikB5SifeQ5Z47nuxKz7iea17JWz8scYnb1Q7NDE55czxBHNmVROC93GEgqt8EdehoGsu3p
fvj3Cm+n40i+6i9CCy+qRC6Rbm9SddOTnuuaHnt3HpEdzTrkvW+IlY8ZSFYDVUkvsLKY1sRkOz/e
mqqU8mwglOEOJBzIjxjtXjK/YSERQ5BbMyrbmFSK+o1SX+n0AbLrBKrmB5wnXVEu+Xi6DinBQMMz
FVVFpVDjMvcycz7Va3U8bhP6IroZ3TwELJJ6kGJDW9xu2Wfm1ZpFxB3QJk83chhZ4L+q1mncuUQw
5exWHyBPfEeEwreiEluImpmNaIU2v7gRx0XxpbdpjjpFDG9zG82ZGqDSnpTm87JdrRTo5LITtl9B
SIwj+D6IJLx6eESODdLvJ+scz/1B8Q63Skhj/X7T8g6Wg8LoZIBySvy7YFjY4XGZ+iEK3vCi+Dnd
IYbxUsPF2hNtI453cY2SZ0dZPuXDATfETONxZ1Oy8UgvHuIepUoyqyQpfKwp3XejuHNeDYEf6CJP
wVt6g4g6+BocsqvXZzpHWjrYJPebNkmCakb66D45e4qj13TlIiXUULKLCLIdof4MVKi6B10q5UyD
MQxXJXXCZCXvSFYl0bdte1tS8Hi8oH2LY8p2kNnBxAe919uWlktzdCSp6gUcapZOCWUqO7W6KOn2
jPEw5JMky51DF+J3OaGR3VduOLQ6ctriwF1u91+muawJcrT+pE5dEf48DxLVr92ZVHA46UdUDnrm
3Km5DTt74QNGbE9ZdhGrP1r/bIVL3hAdHO9nQZ9Jvb+yvGNP5dqpP5vS1jER3K3QKlNA/fCiwV+s
4IcvTqo2Jlpb54X1rYE3CHeKp2HY7Dc59TWz5pyUeW2398oHiBwtcJaObPGCEtOwwgP0A1kr6GGF
lHVsiHOrUEfbOSiC9Uk+WSahplt9g3KBxSdGdLuaf7eur6w1f2mKqYuera12HZ/A6+MdyHPXcdf3
faM0Dne3qzTd/m0u6IkErItnLafJx4XNJjCWj8mCoD+Ll4hBYbJAInAgEZ9A4R6dBT069D80xD5A
KYpLw5bc2fCYWkdEmGg0jN+N2lTtWfsI3J+tZ1SyKyxf8usao1dVtrpCguovcfA88YnWLbIYuFE3
OF20OeSXPbH5LDNjP9j7MuWzNSQ7uC5TGYBHwEWXP+AuEOfbYFUpc64gRZOTqyXG3qSQ/g/N00Av
JOMOiYCZw4VXshWxoBAsniavWoCslU4+Of3JjZ83JyN9Y32QvbmGWWBrALUaYcqllzX7Wh6sYV/0
+zmOUYe1g5Ss70K9ptg=
`protect end_protected
