`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nXFrOJTaws3F+GvsGZmprfn+xnlcej1dPDbqUFGH6M1Nk8b8VbcrkytMCN+3IS+K
cs+76ExkNfCmG46A0VPTR7hu7kgZty+oVHD6CiXoGa/KsxpeL6n7MfgOaetbV/Qy
T8SdGxiiF+IzoDcu11Xy1MBN5KfB3+zPaw2f/b3U+Ug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
FEJoUYCeWE6olu+D/j6MWb3MKXdnOflNTnraUFSd+DilHcDfL4PMWtIA+Am32jRL
z3Qv7cR+Bxtyy9aNEG/tXdOum0KPfilte1EMloW/k5aZbCrkitUbrPy8X8EdCGVS
J+oqMbztFbaN+hb0hVWFv9qf82bQ9qFA7vg7XqcksTBOlzDJU7XqSGyTV/e+o+GI
pIQw1WY8PaPwNb+hOP+X9//Lqf3kcOi/7sPkqHHqShEK7i9vkO9sc3EvnG2vtU30
/kS96sTZJuZuIyjj+IM6vajolHnd+8jZidkKtKZ3RNQ3khbl+f1IZXz69Vvc7jFF
xtlgn1S551wR6TSdi03EQ3tbtSo6SPZ4sZGjIu8phgnC7e7eGdfRtV1rMhGXjFNT
FhUYDmrV98L51wL6aEg548F+DckOO+Gmz1kwHqU0y5FIkt2MtW/M1C3XkEyoVXen
GCRsXMlFvVczntibGs0CXfdxqyL96s3T8A8paylxaXWXN1/R+JKIpEAxAOTjalXy
/hKBIST4AR0AESQWHdd4Ex79cGu0PlWmbqf9cHGvVkvs4bM5NxE3NVn0C6gycWjz
VzhDKg3iXtErapVOAxg0GI6eH3T6sw85+xQ7kd/TgpYbMuki0EoWLfikWd64+BmK
JeRhCUwa4yUKvXbvIup7TOQH766LVkiSShwxH/7zlAZwfkgct7b0NIxKTtS2AzRg
ZXZNASFl7kjQb/Mi5hiK5lFnTp0Yox2tfcWyAT40u7+09rzXKqayq3FJNZZiCdG2
FLt28FPVglmRoLLP/D8/UaCLjSB8NCZa/z23vosrz4vSfwtVfciVuKFTtmpgAdSg
3A7VIoRST+hBzx4XT04QV/3ZZfzwxtOcNGP0gdY1V0lwMWHj4zJQaSsgMvrBYp6a
WydM9L/qCLTCNuTftlM6YMELsxACltezdylau1NE9d7HHCC+ESDIdGJbHFTR9D4M
67wmEZEuGR7Srdx34/duWxe3JvzG3A/HVDXlrFHDysIC05KkDnSvdxB0E8grZBss
fvJefFMgbrv9Wnq0Li1/SwW2Y1hQkx2Lm8j6JteENZ04lAtgDNPIPc6Zfz+yHA4/
GdcIeP3a2nbABedlTF2z0Igi02VEj00hS+WLwOl1XPDlxX1nq84H9yS3FBbclegy
MzOzKkFNiUO2l36yJJpScoXZWE2g7R6Y862+v//d0b6wCH0+QUdP2ejXvAlFmvdD
fJGj3Ox6UTa6qf9qyFe0MXRaxaz9O7MPXARKrOa6nhkKQWLCr5i8U5AUP+vxEYyW
zdT1nXPxX3E3T4/O640xKWR8kvCW720DAx2J7GzgMOwiwzflgrvmGfhfUfR51Hwz
18t2IECHtaN8YdWAR0MV0zrzgD3zwUzLTplMQqfj5OGzcgeGEGC2oLDEEQo6M8GS
f9Mn+NkKTomJU6nnMCvfIOPbyVJskCIhvzGWMn182L245QPFd2cKI4pVhl/vN2Bi
RwDDjLAzVLsZ/ihB7of4fvPfsFDs2VRTrc5sNOqUnU2YpUNBKCrRwrcVP/r0i+DM
a2nWgKLJHQ3y10qZ+3YO3+mGGv2rEu348rg8J71udarmrcbZd+0s/6mTnOR3UPpJ
YNzgmTX/EhoA7thHSoBa1IFvzjeb9becT6+0E51Lvx45lOSLwzMc1gPAKWfPYx8o
CSk1CAVjrGLDePy7jW0tJGnls9/FDEBVNCC+vNBeFi7TDqha+PDRy7zS95HagZVo
NJlK4peYN8BgvjtnDM6A1ILxpGrTRhq0Jh17cYZ5vDUXFWb+83uXJJNqQAkBsBHN
xmH69/JDcJtoe9WYSR83hwzQGVtfsSSKepYLudNV9I8Gs2axbvwjtLBR+igVxzIK
wQyqrrFHHXBNs5MNEbPu3WxbZYkfG6jjdN0hb97nTMLBUw85VKX/FEp6rQWXZyE3
SLOIp27MRPYjOg6pfL0R3Cyu0Kx9SmVic5waeCvSA6faA4A5dgWU0Q1vRoejE6CR
97WYD89rQheIrNPovoKVNOPMXLlKUnMpiB/y/DmTbLUI/TXy3SjGicaGgWescijQ
2oqzCIzewZnRXnRtm+FH3pSBdtR/g3mjbY8KywELfD4+twcDkUmC/p1Mhs0wbisl
5chztLny41X20YpEKETFoDUMP0UA0dSG/zOUdyb2GVnNeLAw7xXNPikvuS+CV4hx
QiVTGu9OunJa5UFr8HpEq9C/WGdBzi3YvKLN1Z2+/w1C4HicmAe+wPXa7zEgtf+a
srBYOhkj5ZnMLJ2v4aF3V5+9PniITV1qplfEdTNGpzB5UoLXvImuHy2GnyBgSvsX
HDMcTr/K07+D0Ofzq2M87gesdCzFzD7zMQ9EsnIccdyLEMBqjsko123u3fYfyEth
IrKnwIFk4Rfw+ypJrSXK69WhJU8vsr3LRzPYDC8Ysfr6+kiapzYQStjqkxwR4J7j
UHbx4YPvEcVEBzDyNryID4kd9odNgDeSF8cmfvEMim4am+FjVpVG3JH8fM0oVELZ
tl9UBpMGuFAsVenrUJTSjD9dnjQkZQKNQyXDdEhmdU+5h/Ct1QlHu9pfrLqsXSZv
fXw/9EDJsIbgbJHdu3oWXZfhb7REc3ZE00aGOw97oP+0oJ1Yyez5XupgxVmc0dmB
NmAG4XIEh5Ank5Oh6wyVQARKPRXFUUU1cfJ5hJUqfGwh4I/BGupbxDG1gphMqoZx
0JU9DLryaOVH6/6YfKQiLYwyQhrFMev2t1Lprfc66jhHGUEHme0g+TK+6f5IHmxa
Kj0rhWvKM+lcsB7kWfZ+lzfA74MAI8uHrz6Vx1WqCEnDFOewrFgk1J9c6nehYzc8
LGhv3giwDWPN21YpGvKhy/sPgbdfueSGXgBpl+pEzdl8WaE+yAf5nEuw65fg2pyK
qoGuj+Hjt7uOJRO/q+UeAy3nv5uH5IY4WGPKrDmj+0xuJrD7utLIF5nfyz/xGpn1
YPbo/Mv8jzRUBQXV0pcrtlc0+MGNQkWzUbaWfV1fUeqMNzwjDKVWknLrJ6WmqhMS
JESxjQrjAKyjFe9WjCBATsfZtj3NDCWk0nHbFJfyJrJJR4UVp0zPNOWujs9bIbgS
q2mXzHXBFmPxOCP6emn3yRtnl0r/gs3J2HfafLY9I7Ols/V1BOXhtO2apy7ICdYz
HESBxmuP/tXYCQvh2CLGwVLJS+vljwPfhRSvohcpefchac13jRlSSnbSakcRge0z
cBzyWurmNeZiqHPna13nR7HKRBA85mZQih4+VuHPt+W+sYN0ougGLfil6Y/85Q+7
afQC+SUW3lby+/+E+ULxycViOx+FIp2+m8wEJvq/KJ0x17x34CMQwpF9NuxH8skO
Svrw9YJPcK8R8oVmOvr+7ofNwQUkxdgP8h4EG9qCEIsMScIO004uGtYULdrEHvAG
OWeatGFpqPWoha3KLsltFXYd0VNxXNhvpn5W9Q4EgCxWZTTRlVFYgkBLSN9q2huq
WuQp4oyFOt+ijWPirqeS99PfPFdjff+H2d4Cw2nOFG3J+vtvcObIxeWJuYanAoRW
6rqSCCTq9MzAueh/PYgJMn+AO8DPCRBd7/ah3DXtDlANKF589wVZvPqC8whdA0i9
LyxI0DG+0lbEWRUfLIvqi/Ve2QRrm6ui9kizfGXVMQS6n6IzHeP+nBmIQetaBldM
Hqt4C1FN+fJZzQzC2Q1sIqckth+Wv/XkqcTwcbJbzi4zob/DY7WYYcIOPrJY7s4g
F/OrYfQqYiDe+FtyWRl8v29iD9OfHMLXwuKWVM+R3ojOgkTDd6PxbLs4YAIgczF8
ELq5O2pDE/r3GK/JJX+7T2dXsZCt7jwd34hP+4b1n0ZUNX/UJBPQFtNQZWqf4MTx
PSl2lVBd+Z2Oq58h0Gt2BPEBbrwGcrjWc8ZR7kanxKyZgqBDpGMd5d9Pb8scjLN9
Pn8UrStwZk7S9Exfp6tZi9oGNzz8Z+GHKJ29bysdQ0AhpBMTkViBt1Dpy1GWZhye
mLfAHvcbtnx2Gtxo/GWd2E/ImcR8xDxTcc1mVSiHkit6Wunc/iDcewb0fTJ+bPdS
nhgX1X1JkOuIwFSkSmZPtwaacptIMa6ZippYIJYQD4ndzIwWtkUWZHlsSWtQMwMV
nJDFhZejsCTnjODZuXfQELe/BDUd7ViAYURlgMhIw+sex3jBA5yyIStwzQaX25bo
AhkxhM5cu1J7Z/mNpVFQNtARNanmgxf5Wajsot8ySkkGrBPchcTVNJ2WsWiXUPOr
NNp8w4MdQpKUgvHu06fVI9EhmLD3bw8PEXhu0yfD1mLEqkUHY/8vowBIiRgQadgl
/HZ7L5KDOadCINujnKAO/yF80KGgs0+NkmYHGx0PvVd3i/Yb/i8EGyilqNBYIY49
t/m94g7Uzwp2UQfGcCz5YViPhSwnXNVREkw3ue2l9eY6YO/uPURXTbBlmp5WLG9D
T4mH293gT7tf/3/mF5sjNGh2+ePDJ+lfFRYmD7IBQX8MyrcLxqWmjZ+2u9MZFmHj
Y+72Lr2TQ4Xeit8sXYN8RKvvc2cYjiArIcGAONIWuH5Ae2LcIKEaiB2y9+swP8wL
3O2gIWlQOy2P/5FxTWSqL0clwihsGbSDsmRgy2S/CkfKIujyJ0JzDmWl5poG9hz1
Oqd90BCyZH1ruMzhnNKPel1dU2jb8LMwP3gao8oHXNxs34wAwP/KnnyBBKxaSiQd
GcOAotrRkhtNdutQuSW06Z+ZSqkgPynIQJtgGptn2lRESho2JwJrcWbG8GWLfZZt
Ez/sCqTmffsrWZJu+g7LS3OQYqcbEwZdsck/6Efr0FSCvtC3X5y5eJq6CRzVyMLq
9NQnobniCDb5vehWXZdyvmCAlrqxmbNmHrewQXXqQIqcPxeoRlQM6tsiRo18vTXa
2OvdVIpg0WtSERwK5veFohgI9AC+njCbNHp4fKePbETCqMitPdKevh97V4NU2iTI
lKWKtUeTb9Td9CTlEXS8fbjcnwJXXtcaF/l6jxgA8eGCYG0ngPS7jJZL+cOhBSpX
FC2VeMW7maA75lTTOfDTuK1BlqKpg0sJ7G2pvTwmVejgs6CY/zIjNdpfCnahscYv
0fDJGIPaCJGnB4xQlYJwhaudjN2hBrNAyZt8b69HE+8l1q38L6gQe1gmlavYpUAP
sCLSwFeTNUmTR9r6Ab086GTId8Mo8i4RGE3v5Ma5E7CGd6dIXUb7d69THUkorpYr
9Rev8Je4TcI3SJ0q+AY08Efsk61Tg+OxeFhzBpwtyKyrKHDI/nI0K2mDFZNcbJS5
WJRZAJXB07w7jHJIZnfKIaTyJK49kMfMsUNpCtG/JPXFoa0aSi1CZBuEifgcd1dU
JxN9x0a66TuWp2MZEXybfsJBfal3ixsXjc3CYvvYicHt8B2dB69Xjn9SRX/xnvNx
BoGMTH2umsdCmjZlj0iSB9bm+J8xiDgQiHydosYrMNQCL7q8dNV0zCaOq5T3AtcD
IoZd0OmobPsMaMZPxl4Pnq/DJClKwwWlQFxB9oZ+Zsj1bzM89t9VO2/HdrJY2f0V
jXiwoJMU+nT2LWiI973TTHdQ1hv+GQWU1GPhv7dj3Cpz+whsk9yS2F3c/VUXv8zd
sQbmqkRzIhEAu0gFmF7wIhU58RroGcROAl7/oDBs9tNraNrUYzo6BKYtUf9b7ZuE
lEOQdILGtMGJGkK69WnY/FpmiodM1aaukSVVfQUSeUrFpkeh8PCQcKsDM16szcDW
Ob+47i+0CWWaER8AJdawA7QRTlJ2ppKxdrv2xwGTbjHDCoNjxW8hOFEBrHtnf/ni
TEUwuFjHWFyWKIOnK5tWe1CbqFIHONvbcaDZxwppkeVdAo7atXVmg5/igZN194EL
qQNgIC78MsGYbqOETdIXC4FUh1AZFL04AvgnUYe98Uw07VHGHLhdFn1KD4qW69Z/
9h0WI9Kt4TFSytbvr9EIVviAeoMht5lyTUHeH6vlLtp9RSNjS5Ajhjaz4LP/bs19
SWkECwrG9oT5GrQCU9HzrSeL1Du0auOb4e1TGsnVAzfxRAC9HZdgndB6wP8RdWWA
IiKROBy0PZUwA2otqp3quLJ+EDaWtfrH9bVBXfqTr4rCDZFumoxHWru/0YrIatuo
foKGGDX5Z2eIgPNSnI8tOhSDsLSfQ8SCEiZY/ikG9U/Ba1UEVnES7cd6N964TE1T
P0Uu/kUA2xOLWUmy9ZlvhjqV+/nlDu/HcIItRi14mRYGEuUnPLPBESrA7W3VJLpt
HHv2/kT6FD6HVqZVTs1UCGrUV1vNqFCAasUjUIkiTw5a0pGZLdYff5IuYilILz3I
LILaa5FU460bBpsqVDL6qzgjerWPpbySXVSiP9melmxh+2+CicBRseCGOM5CnsEB
s/0ZtD3HfGlIHGBS4GmPNn35SbaK9gGJG/0J5HW/tY4g7oMFhE6B+QI7nNXNx3PT
ESCV7sxAAsXEjVY2QNRCTmBVnUHVmiYLUMeWjUEIy9CjsUyAn5K5Mk/e4zbAlsZx
8B1BWS/t5TjPb2ngdU8DQRC+kKG+tj7I5AJOZCNhv+iu7vwi5HuyMkH/InUiYDiN
jgMTKe2Jf7O3IWuAdd1Ea8UPcEqe8Px+ODpynLlv7rW1yC7i7gesJ71+BXxP0H+e
7WPpUgz7CeGR4tNo4s5wCdYXTgSBlTFEiHXHX96deKi0m2HWy8HXz2yXd0cA8IR1
0WN2islUJoKbnEh+XKppD/ds/o/mHxWQaeNc7JRICc8neL3/B278tBA1yGVaSH46
k2ay+M5EXLgU4ZqAHjrAS1S4KWroOclub6gOAzJzuzcvO8TZK+s+jJzCfoVYIp+K
veGrMVpDF1bpPbZAeRCelrVyJKrVvgIsbigL88KyQv9u33EeU823kwNfx6bOM3EF
t1nRhAnLmgXGO0u3BAqAG1bw+9LimXdU9HXeQw6938Ko2ppM2LWxZBNFXMuX1Y4r
csSqOJz4SHNM8L24yCoWuegibHOynC9XJWcYxyJo/OCfUFImrP4dFG68O57j8hV3
UVptz7kGXtoTL6c+BWSe8LCHpBaDrgoYfX/Mqh3QLTfyb9D/Y4xtOVqEmgePKXVr
1Fsjd3fFWwa4IkJxiKh7Lsx/MI1BwSBxUsigm0fvKrFtYaynKPL4lAWHgWh+6V4G
zNiMl3CcRKibToJMdzR5wQS3e5pJTayr2BT+gWmGDseA/ku0lCVkHn3AOk1YFw6u
u+L3F+KvHXu+K9XFz74XKMS6ju64v6HaxJOcnoshWMlAc/6y/GUDZRFcC462UU4i
j2gNw2y+wX9USnuRu3gGPBYA37y4OecxriwJ6IhhKk7vIxmAe0Mtj9E9i/EISa3h
u6WiqLYCGJtYEf7CiI49AKRZgMG+Da9i7+IExv/lzcWPaP83U9sjTTeqsjS/Z1H2
yleMExHQr+yUFneCkehu/Fu9+gLEbdr39Hox7x7W/4KwnSQgp1eLqVaeVfDJT0ap
kRffRauWI0XjD4DCkFjiJ+k0aFjyhjTTtignf2WWgSgdtpkfu+dT+3HZOxdy0mOj
GlEpFO42hTi9OWraVZRXyxg9zIJEPfC873s+d7gssQT7pdFaK3KYZ7wBwganeP5n
JMyf9lvCTHNOglRe/+rRmwcNy3tRrZAIrGmsURWj1zSwV9wU5vIaUuCDCvxWTR4i
db62eq5DvVAnMPtqjqBDwbb1vP6qftmGtrm3pKYRIq+p9/8GINTtRFcoZfeLV+mq
gHreJvFnlU4ShFazuQUqyUHFA2Un4j3PozwQ5dFPvjFSeF3R5VDY6ueutbtv+NSc
D52Mw82grkJQBfp7slqfasPabV+8qquNj+WQ0MosfuFHoDNhLG4KIsLpR3jALcP5
UeFj982KSm2hYxXgpgh9hiVl4sb9fi394q7aSRfZObca6CN9y37T2Dosib5qcFqh
LJur6tu8rFdkTS9XjdBCtwMOcCuXLwx78PzUFuF7JVf1B0lEBUoEXiCXtHx7OqrF
5nq1EOjq7UVLuhIjydBQbgPdsg+BIQ4+05Ie/yJ1twPv1Yqr1rVpnOXKt0gbkv0v
Od7tiZf1qFF+beZclY5fqUHrKrtPpYFCCDEkCz8MNq4oUluZHGPt0/ireJ2mm9vc
QM4NBaguhlQt5s/GlGXLQYF3MEDxHc1JOisin7dio474zUK4gsCu4KMyNPLVQ+AO
0nHSqJ1XYNyPypVaQ/l69Mbu1hdwwbR1r2rfoI+tAPIPYlAVXjSysBgfU1Ch/qyS
WLNLEungjjFQEitQAxz9tbstJa3LoXPqt524jpWtbxs8L35y9CxmFEozN9r7TJKb
sYTtaxh56/IaKgX72I3ValqTFOP19uLGM3TyJY9ZxrEWN3cBJJ1pSJjmhne+oAL4
nBYZwLkKjbRQWaXUnMBy2JDP4lywsHP050uxlDHQCciLyrGNz4Qx+G9GffWBNtsf
LCnac/C1QI1yfhpJtk1uoGzkEzD3O8NHqRnl3DHl5YzXj+c4YlW5Nw0T1QGnq76A
AmjmJsXzyYhwitkQNO2u1SGJMlyQrWxD1b98JPA7vdtNccnhTdtCG9BUNKvSxoUo
qiIW35Q9O3goHvuuB5VXHXQ57w1vw03mNc8q6Fbf9nHKsRJ/uzIKRTpenTOskw9Q
Bu+JTOTgviDD3YEqQJBqY7Gu2OHBZbw2jmjXzimrK5aW2oooUvnJnF9ULJE4GZEy
Hg7Oa6gu9oqS8bNVreKkAl8lncNc+WsraxQ1MWr+dyMxYipdL4zI8sw4ZSt27j/E
J9dHbICW6Ruls4Qp2FLC6SIhFRCGgzSa4aCuJ8THml/jJ+jRfcnV7/i8eoXlf4Ui
MQwujhT+JsUkeAwoY/SkWXehmj6xDAC/LoyBS4mjcpD1RT4JART33yFIdH9wRL4J
zKNt4lqFzSNfyBp32ny7+577f088uyVDU9nftpYzYSJ95WJVV54sxwOz0cAyMcFi
RqpZ3hWCRHFlRR/pHjOoM8njTqyaZi6poLD2ayq7NzJpSVd2sB6H7c+I19bey2Wj
aqCcUnL9szBw2d7jV+Eo7dAazta1fpsIrB+ZeaLTYVFBoppajtEhrfibP4kdAFtr
UhVV+jlQJOfaSkLL6Qe94FjvNLBAK4CXkfkxHw1w+0B7ACtGrEKzMV7ENMH0oFla
CIUN6/OpcoQlNlsGGOaeDP0XDa2YMV3UaLSA4Jg4rsFGVwizdIbJg5I3jbx7KpJe
WPo8lRs9/kOVjR7jNLN79PK9ughM6H7+JOnnd4eg06+HqeArCNwh/R1wuDkCYY+m
6ilpvkWYGS4LEQdQS2kaUeHQ9YYuO6OfhENMCiqkWQRiEpMlueB7F9Quju5pdizv
pVc1jXfJhUTFi9qovM9b01H90zQ7tGZCSWSesRpAJv/a6hq43vypAFH3HSjCGNnW
X7ieYcO38O0rDoOtOeJcS/kRhp4i6/+bCWHpiGMQXwojrEpGQxHeLVKdVtJhbRd3
k/s09k42+cMO8PboVQg1tnKPhq2BSaIh0trMVZtswGi8Qx5LHuz4+r1QDKyKUR+8
eUs3qQsTtprZev4iv6Fz/7FwcZZa68BMtPp4t02Ro7nsXaN4MISO7kTauFvmMlpL
/djNX1z5D5YytBWfIBiB6lLnZDWJGA2afVX4UlHrIJS2sVtV5/Ps8j0G4fW/xChM
hN6Vu/5x+sXMVb6cMy/pDoomk/q3sPpDw+VWtr1172KutfvTIMCGFLA2bnPy92cE
1GsT0zIxh4VeWNv/HvVLhbn3M+JozpQkUvGGpWAZtCZyiDvw5uxY2MipvThkKZiR
EqHQIa3vkr36d/9E7G/g884pR2GMmu7vsT7ik6zSYrdkkBMnb8GHiDIqe7mfEE7H
S8GdnulgBanCbMLdPTO3rj1ny3RcQPTWdSsdcNWIMtBvWEzfikk4DNK07UzIfa2N
qSjiZEBcL1I7EFbAM2CwVLV76EKXTahZgkRuG+WWrYv39m0FgpIzwqE69Ybl1DBr
yENu3/9bnBz208AXl3AaWrVYnbhU+HW9wsC/I7zDUlEDA+aET4yR/CoByr4dK3cU
0rtsZZoj7fOrbfEDfFjlRGZonLqdAwsCtl7UXoFrJ+UQOURP+F0E7s5YfGl8VAli
1xp2zP37n/ySRUerZEarS+9N4HGfz88TLf9kRDGlLXc+xYYx37zk/4Y31AvwBGDq
3O+gEWIiRLBGTxiouW/4K6ED9M2kjg9bZDiEOzGmv6cltbNhR1+GpuErVdf5K1YZ
KnK7IFEmszwWktKx2VKCYp2W1PcGr+6fWqUpwQlokoE9NQXK1MYizVTWVwWJfBSQ
ptQ8qv0Mxc1gj+Gt/OixbUhpDa/ezjibdMaIBD5zI49LvJaK1GbwOIIonx3+Pdjy
XL2IZ/kWfbfebIG8O9yo/h/UftAn3KjSWE9BDc0gej5BCXYgkznUJeDHKkvt9FmP
y68/mPMhjZCuaWbNtkSLfOBSl7ziiBC2v/ZxshARxMKrEpTEFP6JNj0C//U8DiqQ
BAlCBbmMndTuTe+e4/0pR19ArGdT/jTxihLGjGBuwg+KSZPd8/JX2H0SKU1IXLx/
8dKyOjSO4d6kgpI34h64UvacR0TPl2SdOvoQ1tLAkK9u3prP9mcIIqCWP3gwygJu
rTML8/yXvMWI1/pzClSdl2iygaasfWhFvQJmbj4bTwkQBOPwdBSDegeoDCmb8YB6
VmMCILNC06mdGJQP8/1HF6jkbWifRqG8NxqPi6XtC1vSSQ9PrQDMzqX0eJ0vDm2y
wzE/tpFQss5nm12Ez3kntjGmzW1VFWfF9x+NhgvPtNZ0VhtXUeFX2mS6YiXS0tT9
4fDPnqQvKxa3BVxXDycz/dfJg5yLiGcTVupCG6FYAIn6JTuHamb3vCutiSRLy4LL
9xnfkn2JhTbnLYgcZK3V/3SKaCR2iimkBTJ+G44vL1lwox6ns3HdvsvVYzC4qJzJ
C7a1HLn0tMe38KkrNus9vzoadJInqqrEQ4YN1etLuE1Sh/eaSmckrms2InxfpVrj
CdrlUiicZhHG//Et12y8lzpVs4I49PxK5d+MYeQYjhxR/uyR+FYLJ7y784c81J4r
JHY6HM0iPzCBGCubdJKDr0XDDQ0A+OQatRq43Uiwtwtz2SpqI11WqPiKQg87dWNI
/vLrqIJyOBwI1MWsNnO31fk2LDTP8KIiCNe8xmLzB1kqrB4EbLmtccwY7MuLAAd/
ZxT2dQWC1v0ltfvq1Ow8Y1FGO3PQDX2ZAZyOm191ij0apY6XUOGj0NLcaZdEN4RQ
GKs4INAUFu2S+7KCQm1soBasRssyoM4FxT1kZKh7wJ4yjj0rH/eZ3XequGu4Y6yw
xR/OBT7i6lIlExIEMjVZ8SHet0C8WR5FGoZ+gUQPo1vcEyQpcI7wrL5yXGX6EZIa
uV4029G2sO+u91eOS5LwxdG32VjjzTJWIwF93EEAaaR5/EorkCDKrVx+lCO0H2VR
uwpWO/Uf1HqPXRXVdS2Cr6NNs8l1J48WKskQZUWiz4ZnmZYN4qJsZff5+NZ86Jhm
hBJ6VhuO+O7QRkyzkR3HXUuyX7uAyOhBpY6lfmRR8EBRPDmAHL8XjrdIr8UZcgM8
6M3ggVh/4Kb2nVgP3IeX3nCc1PDTFXD3Z8v4G6VbH7bZ9treMeareh7TKO9SKCRH
H3DSuQOzG0vF+5ItFkDRK3n58qcoTDvY2+RXNThOLA4jEIwIF46vjlI8965uGXjz
OQDdbJictH6pA6CvsmpHeJYQ1H5RI2t9vnNJkSsmDEBRAoskfzzTyQ9mnhLi3MHH
sFnh8P5cA2nk6i+JBmT8WUJlmxqu6j9n0gmddAUOz20ARq6swKtCgcDTgRkmdWTD
QJiBuwxA/1pOeLTIxrqdFATU+t0+6yPZpeC2Im6YV7cUI8XfSW8qrBJVnPn0i6Xv
NPqrkafx7Cuv5Ac9SOERxgOP+2cuEI+WYnqn2Cmbuf31g5YBHru2ucjkHZV1tGhR
is1Gsk3XvR+s+pKRhNE6D1RRRw7rHJR/PQLFhOZPMgm04S6ygAjHUi7+S1Hx/3Fp
9TIZ88qBZxgC5zeeyjasMPozDdOWQ8WVlhZ1b6yG954GdY3UEzuUuI4sMmKg5Qzo
04QIQjAkahRXpbIE7LG200G+MAupps/SH0nQIArDvGwfZ9Cgz4gpFo8FywrIQFU2
8FZlPxpTVjyvl49BQ7/IbPxdnnuwUI+CCV4W129CBImAB1yZEZmxt6725Fo5Lg/P
hQ9nyGfADYlhwBNAK/vY6T3xDqxeUVkL/bd9/bEgmQ0I8eQ0nxIh+nt0qKdp3vi8
h8JnPIHFro/l4BGoyGeqFRTZ8ndbhf+PBMPu+lEE5I0bNzPAtRw7bVfszkZqaSkj
Iub4/O9ky/SePbM0jcNQZjMSJMjzzJ46OJz2vTIqzomk6EqJEkvLx5XxEtsZWYkV
kvHxqwmqpU+4sh+bLhLQVTGkaa0EwzvYqH1nMlJ8CSUpkX0HChp54+Wzdsao225y
GDC2Bw8TdzF/5+tJU3I3PbV1XXWqPwQW2XEpXz0dtLn8PQzR3FNuSBYefdlGsjTL
Nd58RdBonpDJ+aiJ0/fTIayEYchNPw9JbF3NxHAtMW9CY39BZRtpEG7kBtpMMHRn
V6gTBzanOwdG5W4y24eSZfy0tdYMuYg7rAqXUexeFbCCyqiqBvgoA0y35hcSlmAI
0OWFAs6TGZBtzdf+i9f91kUe7NZD9klZfy0aIsobvYES7N3RdfNf43Vh77PNOdXV
RTYqbs3OZaXYerlpLMKpxqRDfn6FCSpgmtPfFYPKACMMJ3jEUTzo7oqYXtJfwHE4
1Is+FM71MKR9wpU0/MSdz7kHL9Nnxy2AlTPV9I/kQ+WBqh+uD4PvFHRSWexQy4eA
OYBu3ta7/62cVGyytBc0jSaBI5tv0qSCGtKo15rUfxDGr7iNRlrmA61EI37xO6uy
cEZwlmhg0PbqFB7QQUXq+DyXeBMrB/CdL19BiBYwDWefXwlBdwzPKNQf9NliOp3E
AG+eWBYtl2boqxLwxAdy/jPKW/JY4jXg8p36fGpEQvPDARuFMRJSBPSK9pWUO3WZ
kDdPVjPVRHx/uY4jkoEp5DeZ4Bm/qRvZi8gCGTqpKOd+DPYS5byPVAOm7ZCNBBUr
xi2Nx85pDAllRO/RgkJLNyJtx7JgAQPso2nq9tWTy3nPHf9jCHDJYE12GAAX12j3
ZdUqkh4NFhepH6IZwX2b7ClnnXo8cHArL4E5zgJ/sUCGOIcQn0N37gRmJxrK5jgo
PuLYSdUQeBfXKtEk4XkvHHUzokQq5oUvX5BjVHYrvgyIm0aY5cX5qOQeHH3DobmN
j2KTy4gVvFTXOJ/3mT1mete1D3l17TdVYeqkH7tsc1C54Deux699KsHEp3oDa5XZ
ggdOgKrlCdkPw46BX9Wr7V0ODdaVMCesWE164+i4lwJjpxth5gVBWbIFO6BKFsug
gnkyzodhXpEwGx/icGGavBYvBz+JoXqFXUgR9RmYPPQ3LbVVfXDWdlzbamDQals5
RlXlIsklwETOtpEu3HXW2TSQG7WyT+1WunyOF4Zk2GxdgfvPMpn4vHxdER0bUHY0
St/d++y9koBcPZERw/XWTCmfeKuQC1eCAaAXNhQ0cfk+MSD2QS0RGjp5RBQPE677
s3jIiHFBZiLkvY/4Z2bPSmOHUKcLEr+mUEeuMUnpN4L6i3/ebG/oufQ6dSDx6YQR
rS6C8Hiwe/1hT527uOlRMweR+1DIXi0EKP4xpakm2loN0ZU3nrO93SxRy5TLe6B+
EnPFB6gjGF8vttCVO1r5jo+29nW5ryI3fbo6fSjSi/18hEqyIYE8I899bBC1aKpE
KVpvSlfl3HL2jtcH1Fzi4pPEzfjtSpFPf6H6UB71mi7nitW+61Tw4hb2MpLWnqFU
z1J66IB/TIYxR3jkZvNdPSLV/iJWBiYJUp2EUrhuKAFlEUVQof/GiViQQicDevd7
c1WSBAvM/iC7v87e/j6DCx5pBTr1VnOPiFhE1BbWFdcCGI3SVkkJ3p74KC5YnGMM
8uHCTzvH9l9liGowvbrTnP1Bsamfhq9JIDCxrsmMESF9pK2Rn5lpBrb6NCfLB/0X
BeBjkKE5oiauLdDjq/ESHmlVeEqIYf0Vd23aki0SaaL8fAbJ6ePyrYiKjJV8w1dm
wfOhNsfXB6X0dSwMb9t3oIgNz9ZTpYpVyuZaZfYx+qGeQrpFVf07Wg8bjl/hQiji
vKk3qprHuk/mTgSMbCMHndERkJzFUibONhmcQGR3IkLOG1rxF/rBa/Ec/pHcmQo5
e0hfAlSnxBXcyBTDnMl4/yp9o2GPB557Yw5SiPvr64leh5rpAPz4FejmvCE0LIAO
JIw6frx8F5UJEl+cSqyXbdXAnreCtNZFGcLqMsO6rpDCqutJsu5BHfzQR1Zc4H0a
SlNwHl6esjGB3WwmLcm0hyLN+FLTsU831E/hCGG+mFZi2T0Tjbo4PoEzHOrz6DMT
ElwABd/uz4z2yV5w4asuGuP4eYxMB4+yHKAZrHF+Kcggzf0FANhVkzMzHFeQZGLp
j3pXvgHkDvQp6mxpipfAQcTBnnmGMVi4rfPrDmVRcx25YLcULPiqKzWC6uGf4kij
VOGgLu65RUi96QKWKIGzJ7q1Cc/ODaagh57ncBZXhpK1PhJ8vmCCv9igCsiau+jU
kNiBIrrtjc0oetxnNYP1nQv007eClokydPj8J+/YEDdLozAcy1Lm7hOS06MAz5F4
bUFizwanb3l+7rOGoTeT4xp2ErXXY3t/aiBVP6ZP8EhyAp4Rm86gy4elO49Sxaa8
ifwc6J1rQ6Nhj215AGNLerlh+tTnEnIJJXr7tXDS2thSOOopp/0k3oYUOXosUYyy
4jLJeXBksyUKW/JCgpJhFAI+tgGNAq+f8ia2mNdRz7237GiC7vtYDB9pHNhQYP+Y
5DDx6xiQnHepbtOTdgekygcgQC6cI1JrM9oVzmOE6HSiKPkaP04bOwPQ7mUUB6Hr
n5HfIuE7ZRy2WJ7R6I//Hw==
`pragma protect end_protected
