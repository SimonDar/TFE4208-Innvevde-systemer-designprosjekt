��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U@W~z,r#��qoYy�}nH��(��|�aU�a��t�:�7k� �M�����l�������w�;J������n��+$���q\�H��)R��0h4E��Z�{�\����3��߱f�]A���I�1�-�*�2���NP���Ha-h$:�a���!�,Jځ��Ұf�0�E�FM`���lnK�Bb�iNq$�W��؆=���z~o`����K�6/��_����nB�Shت�Aj���W�p�����B�g�G�Y�zG�9����߼�B�]���Q1�r��0g*lt�<K�zA��7�յ�ش2$7���2{x��1@�[� y���S�Q{�i/� b����2�8\������f8�t�v]ݿu~�7�� ���R?+c��r�;���Y	�;Ea7�f��0)b��'Q�n%�������A�ڬKm��}
����R��$z����~���?��U�r"��Q��_�O���*d���LW�sɡf%��ګ�O ��x�Y�u?�]R����.,ͣU���-�؋�U��߮a^X��V8�$S�B���Ku�8�d�� r�߲��qKl�#'bO_�84X�˼q_Y�ĸ�n�a�22O�d�H�}Õ��.�*�!Ŗ���¹�(BN�F���g|��y,$N!ӬJ}hZ��@�jbm<�*�J��׵~]^�y��[#ڻ�x#�@b��Z��ΰ�p��k��O�:K�5﬎�=;c8@^GB8%����3���0X��>M� ��҇��8���IO��ÂΞ�q�QV_#I9�j�����}��g��x?�ɕ�K�C�hʽ�lCZ��z�B��0��vx��r��� �7�Y.�s!�{>R�\#�*<�6��5j���aH��%� ��w�fsr���xH��J��;;p2���K&��ݲO �s�/1F��F�F&�>��fv��o�*J��o������/�/%z6�0A��@�l���ޅ�p�&��"9gM�@��R0{�p�da�Π�ظ)�(�یù>
����,v�GK�{�����v&H=܄$V7���u�^K�R�<c7��~��A$l�L���0����hto�1��G�(NBU�jjv"�.訞�5Qa)M��1H�#�t�xW����k{��V˦=j�.{>x��ĀG�0�
lf�v[M�%z��0���\�_���a���ݝ��"y��)e�'(e��������ץ�"}t�B<�t�w�8��I4*��j�ݰ`����O�ջfN��ݗ�rum
a�Y�=��	J�����47F3�������
9�跅l�NGQT������Pq�<����48��v@!�ܥ�BӴ�-|Db����)6/t7��B*H�:���ϱ�=��e����gc��v韵��xڟ�R�����4�l�� ��+2,?��>�M��z�p�(���E]��S�-N��PѮ@b��z�DK�߉�JΣ�̿��]f��+�̿��m�O�=M��^s� ��B$B�Qާ���|݅�A4�'Yi�5�6�Zg��>}Yj	����!��I����eD�O�� ����l�M9:����z	%v�/��3��_+��~��x�̈49d�a�䓩��ϡ�^4�K�!�S�g��<����3uK���U��%JQM�_:��Vj�6�}���$����D�`��J[,��2��%�U臰&:��I���o��m��k�J��/�x����0X�?ky뭤���l]0t� d��Ģ�Q�1�̭�^�em����gUj��A�fP�d�4�aD��}sճ #m��}ި\�1�Shq�
[�,뵁%��,����v���r��y|��dh�o��OC��0�F �Wz���Trt"��D����J@I0�1uWBփ�T��j�q�IgS�[*ޭ�:01R�Vk���	7��h�:ˮXkߔ勞׋�)���x^=�E�"{�]jIH��y"�Q/R�k���i�����D��kc�+�݀�	�����:�T6�u��]�)n������bNS�}�ro� ,�ԟ�*vv|��1&��P>cF��"�ڙ�B��V��?�@؆N���W	��V�U)L�$���_ɗO���],�c�����>���Q�k����0yڌ���U��
"���k�0n=#\Ǭ����%�9jR�=΋,�ߗ^2�����ԕd���B4�~�X�
<�Sr�Q?x�&�X�W����v���SY�3���lhǞ����WVo~����!F�N��w�{XjIdVÉ7r�Uu6%�v�`-�O�i�}�Y�x��p�0��D�o�����\�ԕ�ޫeT�����,�A�S�SY���>�@|����Ý���� rZ�jj� ���*��~����V�WS\H�^��ao����������8.�W�ZZ�mȉI�'�g�rk�kO����e���T�2!�Zb(��2��?�ƳHXٜ� -���]�2�U�g^��7��3�j]Q�#I��V�4σ�\��`�=&Ҙ���܈�9�����8��F�N�
��ٺ@�ȶ�-�}�Kv�Ļ�R�ج��@|՘���!�{<�n5���B�w��(��4�z$��;�\k��l~F4�
lǘ��OH#!��;s���蕇�9������������\��,{��8�p����R ��+,4\���D���s�z+���_W(�-�z�� ����]���]/�8#>-iXh�"�U�3�bN��ٟNu���Q>�AƮ��$�W�R�֯u�$�j�5���g}C��vI�/Us�u}�:>��+���[4�|�"��(�d��Y.�G�`?�ԟKy�+�����zFK��ؤ*��p�u�Ʈ�'����y��A�Z�r�~���	g��"[�1��z����<�ډ��'W��V1���x�!p�v�5����2�z�������I�Z�s'w��9��+�:I,�Y�\M�P|G��ס��!0Y4�x���"�t�8����	�e���9X�"�*.��2��i4�c�u�V�c\�(	ĵ�q���@N��Y�ЉZ��VЏ��+���窡�z��x�,wņ�2s}��>B��bߺ���(�����m�*A��.� ���ԉDs]eJc�4�y?-Y�h`�Q}���fvl�b�O"`Z�1��/Q�.�G֮��_pܣ��A���7[��&%_��X��7�!W��I�D����C�9v�{�BO[R�F�5�E7�h������o�������^G1ƾv�� e@?��oz�����@^6T�����#�(��+
�w�$pnQ��,�v�����Ϫ�h�~Ʉ]���Z���$���pxǵ)Υ�ʒe�N[Nʮ�O��5k;<B�uT>�t�幞�u��qd��t���+��j��}29R��s���g+�We@��ª��@��;W���7��)�/H�ت�<����§���`ܣ��xx���*�nT)ź�Q�M����"����e���A.�*!�0���Gp�?���3���?*��mà&��_1�6�
�,Ȩ�9�i	��Z�+�X�g����g����<�@��M�	[�8fw�b(��Ğ��X�M`�l˚@4}�'7̌ȕlYG���5?#�N��4�B�T���Y�v:$�P8s����0c�-J'��?�k� �g��/ד�?�����]�I4�uU4tO�sV�f+��St<T+�5���e�'z?�k&!�|�IAʅ��v��N�Ћ�I��-���:h����Cj�I测�*$mX�?5�2a�x��$G���<�T������GQz-���fK�r��NH�i�H�^�!�S��N�yX���gyr�������c�@%(#V����}����iZ�2Xw2O��nOY��������\V�)1���Ra�T��4�iKF`��W�a��<�%�(�Z�6���A#�`��Z2�0)�H7 �m�)�q��vxY��}r���èr��gr�/u��%8#�\R4�f.�Ҩ��<�*��U����-=��Pf3�GN5?g�bl�A�RD��4�Тuw�%��5a�u��)�|O��,���4�	�3P�G	Og� ٟ0��v:�d��&S�/�U4:1x�B��T�:O����N�KM�%��[hA,���b��[`�M_�O��가B���������:��sNS]���i���f�m��P�j���>?{f��6�G+���v�F��	Gy��8�
�.`��b�/X���{U����y���,j�?Wn����cv	���X�O*q<=3j���e�5x��d]v�̥��?ri���'}�j�&7Լ�iB@��0���>�����S�b1� niqQVV���8����?�I�,�NW����� �j�0}��@��_0�z��}�"�c�8���D6���%�/� +@�%^�#{��X��=��h#��r�J�(�-��:�\P������vg��P���� �I�IU��Q�Z(����W/2���kh�Zf����-�D<�r�(��Kә��*3-��-�z�j��yJ�}���tQ	��I\*{�u-x���^՜�rLwf��;�h]UH�̱��("GB<Ox2u{����8�gX�s%"���m$���d��:� Q5V�lyx�^��As��]Ҭ+�_�g�%U��%�Àq�=�G�f�{ǜ�D�@'���ıqU�.ߛ�WiF t @�dEs����E�g}�p�`%�̈��},0��d��R�Qɸ�-�uR ��m-�-+�3
��q'�X�C 8�g��LG�0Y��z������P�4Mus�dm?�բݟ�b?z��Ȯ�cr����Ҵġ~�>B��A�ݕ�ރT+��sK$͑��qT�V?8;6�)O���c�/r�H c�庣�YK9����5뇿���]��_��ҳ�q�²�;�PS�Rt�N���g����A�d!3��1:pX�� ,G��B^K1΋F�bk�g	pC���A%!��A>�o��p�)���oy��O V�i?h,EZz����"�+]�4��y�+�s4�H�}���!7�$Xv�����\'8���}�bzlve�!�FD�5[�2��HYtv��4��0*�K�V��@�-=��ش����56��<�$v��  ��c�+��	�6��Pe�3mF{e�f�V�����Nn"����¼���VS�{�#{�&>�f�' �e���	o�+d�[p�_�{@T�7|�����os�������k"o ��+:���|O�(M*�p���1��k��*��qn507"�ʎ_7���p��xi?�16���7F,���c�.ކ�j% �(OaN���CwW�i���az|��
k3��<d:���՗��k<Q'%S7]��c�LF��v��m����wԱ�E�xNI�݁V��Rn��*�����94ʅ@�Չ�3:CRv��;3~�&7և z���z�"�|�~Ɍ���-���^X�&H��
��4��EG�S����m��Yi�`�k)IIbh��T̬�ՠӁ�0AT߅(^w�:*	��iV��w�<nH��D��\`�����/��]Ŗ�����v������c�?��WҪ��kG��I��o��hp��x��GM�ugcB3���UHi�G"�k���V�%u�]���
{������P7�o>�%��=G���M�`3S�O�Ε?���^��z�]�K�l"n�_ڈ�S�A��KG5w�6��x]��Z�y*��	�9�m�H]IW6���C��t`�1��3<	,�l��RF���	��ŕ�MV�?(�n�{t#�s���t��łFd.1���
N�6k������c�	Њ��f3�Y5 �7a�Zz`���9e�S�Z��;7��lt�s�w�?��I����yR�Ca˫�+��|R7ΤN�2���:ꢷU�&QL�CTpOb�q�6d�H}
r����R���̲x��!iK�c�[�z/���D��ɳ��Y�_-� #��B��%���M��M<������5|'p�4޻�9�o�SB��eN7��$H,z
 ;6��_�N�r�=�� ��_vR,���&&?����YGo�_�y��@�DC=e�bv&�'���T:��XxI����K?&&�),�!��p�ކRh���X��?ܡ�i	>dо�D)�K��ք�!�U�1�w��6��>�Є{z�L�4}��Ņ�����b�I�9���	j�'��� X/���H�P�%h�L������f��-�� ��]�-���z�21��G�o3���[�F���4�X��R�"�f��:Ͼ��e�(�+Q��D���!mv� ����H/T"|r� �\oGS(�(NXP���bƫl�c_��J�_���T�6w'�"��\��ۼ�-������� �r	e()x)P���i��B�RL�}R�jN�$�A=%�h�:<�D9���_���f��.[��u�G��½�4��E�{'l��l8�����UqK�h�� �	�
A�'Xx��_
ꖖI�z:�t�'�(>ڀR�5�NRW�G�T�7�ٖܣC	�&����A�r������-w$;�}�]�Q�c�EJ��3e\ٯ�
�E����ը�J{�\��eW�	d�%����S� �vݚ�1�C�"yQ�����_v�����P+a��I��)�!h~�Rj>o��#f������Cxn/	��k/>,�|(�sz4��i�b�E�~���qfbEyJ�bE���XBLw%�t�w�e!g��M#�
��uq�z�#ؙ�V���Iǹ�_P�0^^^u T=�I�T��Gi�\x�JSi�VtM�h�{���Q��#��9�
r��5����,�Q�yG�X�b�Z�jf��̲�}߉㭹��j��<g���K$~0��Ո��A�'<N�o��NL�܎��;>�aZ.��_6�y�V� �ZN��ۧv42�~��Y&�5�J����й�Î����Ve��XGm��Vwη*?Fq�̥����Ь#�P��n��nɞ����<��j�D@%q7ݶﲫf�(썞��3�������zޮ�����{ �ͻ"���}RM���0;���*]{��d"��(&8��Ks�!6%�?�זJ��A����2]�oY)ҩ��
�;�w��Arf�{�+����5.���ۼ3�IhOŠ�D�������K	��c2dj�ݬ���t��j[�Ґ�f=���E��Sg���9��? ��>��c�5&�����O�C�,[�f�r+ZpH��~��i�D4�C�����l��`ˬqjy�&@q�������Ck턳�k�U��Z��E�+�;ŁtyGp�+#|3o�g��O��I�;�R��J��Fn��{��!���\n��"���	P��'s�Ɇ���B�1��x�zū�c�w6 �md� 3Q�gC�b�>Je88c&�h��Y����At6t�]��!��Ʋ��D`#|'��EdX��G.�׿����������/@dY�n2�T���-��a�'Q�
��/�@����q��l��3@чj���;j8��>+zds�q�s�վ��.)N0��;�u�N�FݼO��x˧�ܝ8Y��J�9HM��TтY��÷#��囜��0���B_��-kEX�$���E8ؐ�= �T�:<\o�A_�o�Ѩ�P.�JҚ�J��!<��&���x�%������Z�����ޕ�l���o�.���}��D��簧!ч��H���!ܝ׵&?H[�Z5�-M�N0Wn:�8֊�{"�5R!��j�P@�Y�Be|*�J@��wXQ���sD��'��a@/��N�6r]EV#�+�I��[�(�;P�=cX�@�?�֬����$��Y����s���	u�=�4s/ׂqb�s(	�,��@(�Z7�PD�'9�D�VUV�9R)
���U:/�si?�s�D$���*X���k��Ča�M�������DZ������� U�ф�:� [�����dX"K�&�����A�aM�����[��fmb�k�<X隽��[�o�)���~,L	@��ه"�sNG�ڰ��I��� �X��<��g�N�&�?53аEŌ���z��!�����[���%�H]�~��*��4����=��6��pr�j���5O���N���XOn$T
Q�aA]�i%`�lM��e_K�̌�Zq��m9� ��ɑ/�yf�2�5Y�^�<�Պkє<�Y��6\-�161CJΆ�'_�N.�.�����1����Y�X���/c�ڇ�D$�p��\�y�[�����!�
y�6���ͯ�j8��~o�B���~��y���V)�N�-���2]����J[M�o.k��,���o��s�ڇ�1�Y����� ���9V���p�:	���G�;�r1z%I�Eԟv�Z�<�o����g��p�,4F޽��b�Ȳ���Z}�>_`�~![�<W<��`�JXq�E֜�a�}g�L+���t��4��ExZ��\.m���s��ym-lT��T�!ͱ�!��
�X+�GR�%����&Ǽ}�Z.�F�ǩf��6�='��Dd�dO�P�τ�O~��b�W��^��k�|�n,�>+�ƻ���)C�We�Yhֽ��:�(������[v�h�i��Ǟk��8D凴�_�����[yj�ڠ��c�X�_-�����������Z��q���X�}Un6��(��&
���ʥF�jE˅ө;(hgD�8�Űv��ߓ�����N�����j=x�1UY2Bvo�|~:��zy丕Q�i�m7x+�ϊ���	�"�l��Nj��'
~ΡpQ�:�[�"�t�k`�~翩	��&.9E�B6.+&��Zf1�0t�0�t�+�2Н/e����r�\"I�n�>`[p����@�>�� ��X��vϒ��D���Y�D�kT�-ק%��o�B�d̒ 㽒Բwu�9�B�m��� <~�.���T H�N�>F�9�X!��#�H[������#�1�]A�����h�0�^����SH�����O�:�7�g�,�)�%���P�	��o�{XHb�\�����\�m���/�R`i���H#�5Ec8���h��Te*1)�^�����]o��u0ap�`nc��=l�ť�)�Ȇմ��Gx3�s����
	8@���B���h�	��Z��4�����(�����M䖿9������S��_�ڀnKvO���h� ��9�d��g �)4���:E@HyMM����i/D�������l9�9<���b��+U�\갋#���xv����}i�mB[�	�����x�|[�B��|<9/!�.�x�*��!��v�|����o��Ť�f^톐ud\-g�^�-�hwA�/���k&�
X��%�X�T�?��/���sI��_���0e���
�~�����}~'X����}�}�x�M�c��f�^RY'1�F[��>m4OѠb����{�Y_�Lא ���A�8�1.̈w<ŵ�����t�E���sx�B?l���m\�_.��k>!��ES=TVh_o�ϑg��?�/_|����P"��ޟ���hG.G�Ol�I`P1��c���'J�%�pZ���]j�"`�ӧ�O������� �s� bf���������g�Іh	���f�940�@oo�aQ�y�����ooB$�S����n�={���2%l�bp�aU�mL�}�:���B��b���DR���?n,C��Pu�*�U���ٲWQ�*�Ʊ��+!'��ɽ�W�Y��H��.�����f޳����Ƣ���3��;_��sg���T��`fO�ڏ�=5G&E6���w��<��Iש�8'�\U�!�b��C���s�X�J�|�X��(��|A����ib6-5s��J6\��.����+pX�.��EdaM�c��%�e4�Tr��C� e6�즗6���AnmO��Ԇ����4���\��|B�DR{��ǫK��e�.�6.�d�Z<>�|t��!���V��m�4l��[�'tH�T(��9p��9r�� �us��₧õ2�3]<?���!	Z8)4�T{͐���SYV )1�RB;R��ni�^ z\d�7J��
�}*���:��5���`�2�Ѷw��A|2�%�v=��.r!��iצ�� 䟕��Z�|�7��H�W���\5�x�1�f�}�ZVa��E5�ş���k��$d?	dmμϘ2�6��q��m#eBV��/pڻ�|NA�+A:������cF�_"A�,�wO���鍀%g���W��O]7;K�� ���%���$��7#�F'�{��@���'K�E�t���QE��ND��jM��\�� �����+jn�I��ƌ+�2�G�pLݟ��_S6��h���H����*S�C�bƐ:���l�=)�[����Z�C8�߮�����-�?BJb��e丸]ev���_]ɨq���[THo��\�V:O��t�,�� 5��9�8�Ao2��mr�k��"�z���uB�E�Q��2+��V�'G�I���<������S�,H_RP)10���ix�_�y���U������W�f-���a,
�\��o �sS�Rb��]ŏ(��\�0{iu�����)A���y�#'����ŝ~��z9���`�h2�����4�u� R�Wc��O�* �@����ĉ�%�JX����KBg���x�Q��6�W����z)G�;���=yYC���+Y�N��dR�34�s�����_뗹�~F�L���\��z��/���T&��G��{��I���^?�c���}�!H������ %��_	Al@$5���J����3���:%x��pM�0�p���
��t�h�����KG�Q����A��j�L�{u���b�u���k��<�Zg֞ÿro�k��0��:]xj��º�NK�"�5N-�f~��y^�8�ӲA-�8������⼽�-����k�B=�WV���GmGDr�K�u	˯�hd����_�Q�����,k�h��GlPVL��ٍ68̩��Jkd�V�x���1�YN�;3��{��ֳWW;�sq� k�J�6����鱧�_'|�o� N������^�|a��D��7q��j�}�0Ȯ���1#�O����K�jo,����:k��q表ddUEL��B[7�Fo������	�����I�Opqr����>4�^C���s%@fV�܄�����3����Yʫ�����o[�:]͑����;��� X2��]��,g�v�9v��q�O�b�Τ��p�O,�^�W1���V~��V1J7gi�C��w��������w;�	�@�D�[�DڎD�M]�xQذ��#��'���Wݣ��Y��5H5�
�����@q9�̃QΛF�����.��e���q������+O���БLo��aB��Bz2����N�H����IVC�8���?9�3�'�W��"�Z�fj��W�e�򏁮�dt��"�Ƥ+�X�B����3^(Ťa<��䔃f^Y�]�+�і�l�<`8v�`��g�0Rx*�Q�ui���'��
�ST����c���&�;���?�h���/f�ܔ��k��ɫ�\d� �>9��`�ۮ>�rg[O�j�1��P
�&�I�������	y�v�%]#��O���o>�m�Z�"��jy6���e������V;a�,�S�@����>���t�7�/� ��I�Y��D$9U��6!Sh�1{�)Oi��O��Э��JU�P?{Y�?��|��G� ��`�P���
�ή�ux����e�v�g�ԫ�2�XT�O���,Bh�d�]D���VPg�p�/��>�;� �A��m���G-{��ױǂ�؇N�-��+�����Wd�$.�KnŬ	����r��="�x�t/�����8��[7~p���D�;�w~X���Z���p�b��=���N��c�#]� �i;������_�ùw@����l����D�f�x\�@-d|����0��XC��5�:��J�P��*���3���.7QtQ�w>�MaO:J�X�ܞa�.C�����]�̤�$�z ��y�^���сѐ�^��,����]�V��zKᢺ�Q9 O�qx���h�ǲ&�� >~��a��l^���ؾ�b)�yWt�f�kO�}���1h�� �i�"X���q�A�E�}�)8bJ`�n)���k��'#��IȻJ���#�#Ր�f��C���v 5��~�!����>�b����ms$�������d�R��`�.8ޔ�D(����)z�ɳ�M��	��.�'�1�W�&�z����+O��+����%=��;6���zs�$�`�6r8~���e� b�82-��>k[��w����� �3V���ǧ��
�o�(������d� ��ބ���o�ks0ȓ�S�x��qc�5��󪯦&`�
��!�W~cn[t.�`/s���\��?Uw�X�i�O5�FE�E��M��f+@s��ڞ�U��%\3>�Hݻ�SS�k�R�MN���Ǽ�X��F�Ɖ��/iڮ{'y��`! ���ht��r�R����u!�c�k
oʛ�<�wxU=Y`����kơ����n����C�k�,��G#����E�;�
�#���(<���_��>��6+�"�D�A:soLxJI(���C�`�%Q�f e�?끘,FF��03M
�^���`�55V�g��ni�!��k�A@(�yAԢ�(Rg����t���b(a�)�v��d_=�&hH�=��鳰z7j|p)h��ss&�H��&�g?^e�5\-�$�\>\@W59���8t_l������P[W�9��t~-qv��(7%4�Y�w8cǰ�sק>�U�E|R���i ~���԰怔�6l�<;]�G�o��찂��\H^��S�i���J����ծ���Q�|��g0�C�iʞHK��L��3���5��#	�%����v �T慷�U�� �~�d��|͜*����oڼ��mZ�Iu#�a\*��P�S��zd��nJ��������ϳ�*�����j	��
a,�g3���RD��oi�O �9����> ��*�.�D���<����&=���c�7�B-x�-���Ϩ3��	ϓ��1�K0�4��6�^�$�� ���:�V+���Yz��M�5֒J#^��+GT��� ў�>�̍-����&D ��yc�B�����q��U�|����AO�HG��h	��+.JLMױ����D���4*S��-�g̗N�Gz�9�!����0ϖ��l����l4����Ͻ�#���D,�}� ��7ַH��Tp$	���l���FK(l�h#�i�ʟ�ˀ-�_�O�(P��r���ܲ�u�f��#*��c�Vry�k��vȩj7�q)�旽��8��!<p�R���o+�+������`�E�z�n��	�KJ�ԜN��q�R�5�?լ!\j2dJ5E�4>�\�Xk�%�*����|]5㶂���0�%����/	n�oԨ�:�gQy4�В����f$����d�T��*��;���!��yu�f�h5Y\ukD�\i��Vd������O��тO��7_��w7#
v��S�{�ޗ������IY#�4!+���W$+3E{��]@�yzK�ձ�M$�Q���G�����1|7y�{?���[�Ջ�^�(P̘�~��,{$W�rr����.�-^E� �^��*z!�4mFA諨��7�W{�n�ıv}��>\�Ag��\�A������oB��՝)��q]�B�a;�^t^�&^��c����C�����Ծ�]�����:� ����]dfH�?��[��A���vrS�맕�e��-ۉ^�P*G=��4�͊~� T��]la>7Ji-b92/膛�pL��F��&@�&Fk�[N���KU@*�cm(�.�X��l��/.k�n��X)A ��R���ԅ
%�â�0�*�7�QX����q���Z���l���ן�V����bB���ꮕs���c{)_�.�3���W�n�q�	��E0�u��MK]Dc"�V�����R�ؚA���Zi °PB沛��-��4���S53,q׳娖F�[C�b�:Ś����r~��3������@ؼ�m��UK�_��Ox'�7ZsN�� J҈�<�*G$F�U�;S��y��=Dێ����op��a���rW��C9t��w�����#2U�#�#�+a��f3�d�t�t�5�ᥲޣw�"����O��%���;Bu���-$H��^��ǆ��M�h�~mH�!�g�q��K�8�,��u���S��âmB���ܫl5��!��͘6  u�G)��R �+EM@U����=.�R{e��.*OfuP�8�������y���Rإ�:�X�;S��]��Ů0�h���ж[�ea�|�����o�n�3J�M�%qӞ����T`��#x�����E���D�X䔻$��M\M��&]pU�e�s^
l�y�s�֚ѕ3��A��Ȯ�Mt)��F���*��)|�S����H��z���<[�~�7qX�<�TNuz���8����O��_e��W�U�<�l�s�����M0x��C��~A���ԝ�N2� ����B-Hi膨?fnX*�U2���6�e�#��T@�v��'4�|� �(U� ���X?�^CU`�|iߪk�|b�p����5 �&X��X�	{�|��c��������h��D��6g):����Qo��p�-;���7��C5;\��u��c-3k�M�&Á���=\Mj?#2ՃnS~�1�Ѓ��V�p��Q��UC n�*�l���L8y#�7}/9��ѳ!`+z�z��@�����k`��`<B�4�ͩ�'��xV*e}���������cS@��:��dP�����PE��M�m�Gz�X��.��[#�i�|��_�~�?e��p�щ���q/��_��y���B�[������`�XΞ4�����S. �5�3��3��ܙ\�M�e⡒���+}��smT���-��v(�D3���|�B"[G�8�8nP>�c��|!Ml��l�6�OB+��
4¬.�:ݒ���wBP#�:e�D��EՆ��$lym~�8[�	ǂφ8 I���Xp�n4���Q�:�k��=�h.{E��'^~0��r5zZ򈺭�/ λ�U\o�Q (��e;�ރ	܂\%	݈����.^~
��N_��^���g-K-��eh�:j��k���n�>6ʋ�c?�1$�kK�6����6Q�1x![v��熯���hR_�+q���`\{����wZc���,C�Ёn�>F"�G,��N��hi��؏Ã�v�.��ZoZ�q^d�2-獎��ա�qfڥ��t�j	�m%�/�R"��$V�}$x��vq�Z�&Mf�Т���_�*��r���1�7�t�$�M+)-H���D����G ��uТ��'�)�u�V�p�p"���d�]�� 7mE$��fBsXW�AO7H~>�P�k�N�̄�KzF�;�~��E�5FF��7�~#=+�$}]p�2����.6��5$���HN�ņQ
wji�y®ˑW`ll>�7�=ˇ 9�&��g=+����!@qy�������u�(�'�-���A�'#�/ y֪��y�ў�2P�h[w��Z`lG$u�q}��֖>� ��A�+�f7��n�F��<d-I��{dT"���7���m ﴂ-� ʼD�x/m�מ��Qv�e��(k�9c�s���>��	����1c�1�mn���~[��`ks�A�&!��� NPN[(H�u��q��|���f��}�o�Q�W𿄻V�������b�}Y� ��).�aޭ�~��`d��:�R}�����NyZĮ�V�������*\b�o@���""e�G�W���R�-��-�d�5��p��j9/����c� 54A�ckct}����^Ii!95�i'����:��:A�,x��݊��1a�*�6c��ZK��� Cp�vo��\�����3��R�N`�L�N�i!��2L���<��D��v���V0�w�����P�K�klz���GcD�I#�{��ġ�8�%r?��.��r�?x�c��6��v���c$���i�γ�h�C���}�1��ܙ�w���6f>p��0�����+{��#�%-���֊�ԑ0e|Ԑ�"
Pj�S�������E�U6!���?��)
Q�͵���qu0}�l��&����g�<��������wWґ���Z�������W�^!!,ŏh��6�֍�_��Æ�b��v�oL���R�Ԁ�fN�`�����Ow�]���Q�]� ^��Z�*�V �w4!%� z�Ɉ�k������D�j��nɶ��iȥɶ���VN	��%�v�ڣZ��Tt���\P�iQ����f�<ԅt̂�H
R�>5p�{�k0�ʍ'��7 N����oB��w��m�x��U���]̀�\N�{�>f6TJ��k(�
ba�IM\�5qA/����C�,%I�������fq��*t�DM�_����C�GC����lN���w��S*B�p�Td��۴9B�����7Es 3�aGI���@��{^_���dDtâj��Z��^��dF	�\WQi,���+�*U�+���`wc�b��qT�b'FV��n	l�K��E���H��>d�^�+�~	�1k��`[��If7����q�\���#����jV��0�~��!�d�S�`�"u�B��ٟ{�[J2͐�s��h�-�T\xZM�{ �QW�a>	�.�����7�عmC�?�V�98��#���D�	lx"�da��N2��ݴ4J������617/�Ԁ򾡲j$��Ax��E�eQ�2N��˰��R���g�����d�����((��o�5�	Һ��(����� ��֨�z���Q��Y*������c`�)�<�`�n@�]�4���-��ĭ��i��!W�x���Jy|K[?��:�����NP�<�ÅD��(�;(���}zY��Re��ʴ$��B� �6Ylq
	�[_~���릣��}��P����;�}5Z�ͦ��7�Ȇm�)�fϾ�ۑb�ɍw@RJa���0��nv���ߦ���R��(O�	4@� ���xzJ�P߫티�J���m�z�&u����k>>���&Е �������#Z�X{�z,B�4>*zz��:�F&��mf��WZ�Ͼ�X3��t.H�'	��H'4�'AH�&�x�?Ĵt�N�Ҳ�N)z���T*FN�z�Q���a�~K5��v�|L�?_���H陥jCN��a�6�J�J�ɇ!w�d��!'����K$/��@��Z`Yr�Cq�#z����TFfHSLqg�M�����ւ<��;�F�D �iV�?�;I
�@�f��$�a*^����K�n��
����rpP���-�l�2���-�O&��e5���9�b�J�ai�U�Q40b����Ad&�b.1��;X ���]�16˶Z*!c�D!�������$���J���.y\T�@�|�0���=$�>;~�*�����Gp`Bn��+��wf��i�<�ױ��[Э�$�{-�_�O?���hu
3A+W�x�_�i1����H��Mi�g���*�=}����
�!���T��^ٝ-������g��0��Nf�����Y���q�����y�͊
��1B*�7Nx�w`p2��`xsK����3<�ꄨ��7�j �c�{HA%�nm��}|�9���0R�8�zxm�G�]���0��O�HX����)��a�^G����7����x��ƙ �o����E��d��\�SO�gi������~K|L,+[����r����/]h;}ǝ�����k�61 ҥ���)R�7\�+�2�u���F��}�S��
��$�Ͼ މf�A�0¹�u�`ߊ�ScȸmR�Z&P|()��>�w�Y�m�_5)�_��8��I*����Ll�Q3��L�P֐J��.ܼv�_E�~�w�@�����6+���>�|
�4��?�Ir%�P���N~�>X��2i����nm>�S���(�R�U���Lm��
�(W��90KZK���ǳ��
.�Gd����E�����&R�i�!���*l��ԣV6���Jf ������Sӛ��a�z!�E�f�%����`���O�L�e_���E�;Q�O�a�?�!�$6��tp����"���F��Џ�&&Sm��eN\h�hEX���C�w��gk`RuJ�W�Ʃ#p��|��W��LO���q3/7��1�]�Uw���w�$f�����v|��T6�D�A��h{��!��M�ܛ�C�	����k��il��6����.�.�_�[V��C�`m��I�*�����F�޾j� N�\��h��%��ܓ0T��K��!���g����S�#^�
tuu�T�إ�,4G�mt�� �{/Hf �M���.믉���2��թ:��ܡ��X}���J�#��Se�<*�e��g�=ץ�vc]��y�:J�%��"��(�:'�r����Nᅂ7>�qJP��4D��	2������);�L~��o܁�BO=���U�4R[�{	 5�@I"�o�c�mKI���O;q���1�f�5�o3��Z�W5�����;���IzK�Qˠ�@XӃ�؅�x�s	皊�^*����C;T��������j7^Z9��B+�d�,�T�ĭ��l��i��|&޴�d^���H�q���`MLl�'�4�e9�������8�z1�r�����&d�7nT5d�a㺓��|�����2��vw��z��nR��_�.��wTN�IpoUמ�v�]�D��#�ߴ���G`��gSw-rbh�K�����ܮ@]��y|�[��J��ek1��"���A�c?�2��3��N)uD�U���].�s�-�� �GlEhάz4�A�/8\l_��|+�i	o!
Z$[V���QD���|�}!�s�U���N�;�h��ߟ0[��b��@��a"�����7�/�����|�<����Ozy�Zj�
����V���ɴ8�@(\+<�8L��ά��h|��j~�(�LZ�������א��V����7����iĐk�~ʓ�M��>:��f�n4����]P�4�c�~ה�ӏ^����U!�"T�}�"'��??J��j=��G�#���[�M���ʺ]�3�/[��Cت�����([������픛k�Z�E-4n�:�� �NŦ�g��S��5��ń��2W�*���6��b��C������P�r��#;��<�b�4��B���b�
������,��$�/z�n�U,����=!�#�'�f������E�<.+	�X�9G�� O�Yoq�l���y;I:�
6��4�r��3��ҳ�%=S��ʯ]e�,��I�w+DX�=J.�B�D�dw�);�pc����yV迗ӊ��U%�� AC���#��8�܏1Ϩ�ͱ���cK�k�T��R��2Grt�ߞ�'�xh(-�7CC�rӯυf������U��ܬćY�����+�����.ių>���˓�Oc���C��7��)��躾�d�2�N�r�U���{M�!uV�����mgY%E�I�2�=J��^�E��%��zn�D���´zhD FF�@t<�!�:�ӞN���� :>|������+}&��O#����398͜��V��zo���-&����:q�vr���/���<�=Ka����R�,F�N�j�����ȴ�?u�z�$H?]��og疋�lG����\�Y�UA{3�kD=&^�gԨ��kXO&3�0�i{
a4��)�߭SB̙��pȷ���(�SR���"��4ݝ�Y�` ���x�M}7��̑�����zֳm�{�KR���r"--��E�9Q���+�/�����˞��E�6�LNܑ���l��G�	?ifsW<Fn]�b��pO��EC��~�ʹ�^{�Z�/0�����	�D�OK�P�<:�p�[f��Y���&'qO������Q"�~
��.�O�y=��d,�����L��/s3���
�V�_�h��t7^��qB��|��0��U�t(��G[�SxE��@ll[�����N/��Rhr|�q�o5 �c�9���E]ޢ���S�r�\�foP�4?�ܬ_Ps����?PqO�]_��������dPV "46F�Q�2��YM���!7��v�qQ�a�6����ueq�l�&���'W�������Lh�\�N��-��uD�X+�H���ٍa�������۬��jb�����rۤk ����ܯ/�� �\-=��_~�ϋG놐�]�A�!n�.H��c��DR���kSշ\���t;(�b�Z��DD��}����'��?��]�a��鄮;��1e�R����^&qT��_�h�j�Hb��{w�E�ClBF����0R��C��H�`i�tX���"UE�#�>�J�gЮ"��t���?�M��K�J]��\"9���3�<o�1D���?aR�$��q�N9��d��jmE1}�.��,7���"�)��H:	l��s�T,�?8@?�p���K�g.y��/R�B⚅!e�f(����ke���QH�z��y��<m�SqX���f�
_[�(#�W�Q�T�b�T ;��L��^!e+(��VӞ��HS`��$�h����r�j;@A�V_�4@��;m,~#Ⱥ��&̋=P�6�2�duc_��(��F2����8���� T�l��� T��X�B�Y�'	�7��<������r3�G�aI�����ޟZ&��!!~�Cl��.%�O�Gw��� ���G�\ �r��9�=TM��i�<���g�[�¹7�7 �u��$p�D��o�C�ًs�k�/4;��u����+�yQS�[6^_ai���YmH��;�)����ou��Q�0/ ������}O�n�i����C`�S���J��0v��_t�����G��^��Zp
��G7�϶�2���)8���^1� 9�-�:Q����$Y�,�~���]�rrƃqtQ���R��Y�n�0����s�#�4�� �e�kM/�}iQ��˟^���2]F��b��㼡�Y���T�P��I'��PM�����YC��?-�-��\K��		�w��ᗞ�0����&eOZ�^���RE�4������qx�P����}t�}պ���pVu3�G�͍駄Q(~6�,8:]�F�О��ƂT!Z�34��3�/�~�x��+A#��fw�=�������72��h)�Ӕ7#�����F����_�մ�3i5��}@��ՠ�p�� k��z=45���H�no�	�%%��Av�@�>��w�)���8�}`�H��j�Fiέ�P��A��F:k" ��_��Ҵ�{�����8�)ٽ��������^�X�'���B��4��b�i�����m�e�p����0��͌�/�e�R;�V)hl�w��W��e!��|�>d77�����q;�M͹d�k�h|CxK��
��9�.���&�����WJ�X�]�xu,\gf�*��!$c&����c�;л�MC�\^@ZiP�~��B�NR�2:�#�Lt���q����������B�FJ��������I���Zd�H�4���잔6F�����%��pL����E�Yj�ʯou����P7'�[m����;OU�$�E��+��t�l�՞0���̉}GԔ�Z�8e���b�~L�,m����ɩ�������I����"�*�rpFZ~�W|Y*��[��T𵻏~əD��lsV8�@_�����<)+��K��KTW�3�e~���G�=bk� 1N���S�>�P�~Qf�a���j���F�/�_�}=���2YS����L����|��*a�T\[�	"���j���Ŕ����ePmu�$��4���_8��C��w��yFށ�j�/���:�i #�@��u�<����z�f�����3<#��V�Ȏ˹%O�$�4�����"3zf���S
�Ɂ�.�'���2�����Hi�0��{&p�e7��&� �+[�g�Q`��0����>�N(�B��=\<ȯ�5�1��f�0+�$��X����-O&��JX���!|��dl��;#LT�r{��UE�~�[Z�f��T�NO^g�����'�P��}��Q�i���_�2ݖob�O������$%����T�d�ZMȚ6�TF�T���*~d^�~�V�?����E(��|Y��N��f�<~y��։TgR;9�x2ڙ�%�*��o`ǋ�o(��P�D��Ϻ����R���6�,ߤ��J��*����d�����C��a"��OM ��T�gy=za ���a1I����)�i�������Kt�<�n� �g���\�<n`m���8����.1}��s�V�>�%���d��S�������N��� �T��\!�+c3��h����,�M���*nX���#{T�OL���s����{?#B��E�ɾ��#=���g\���i���TT`�eG]����˛xh}�/���Icu��Kf��hf����4��M@�����l���i?^疅�J�?���>�!�)q`��o�M������m�]��B�A��7ϊ�PW�e]?K�nY_����.�|`§�/i���Y�A�T5�₟�ȿ=lҾ���H�x��}ҽ���/��۽�y�Ϣ�lh�ʦ6\9���I��30k?�d�'N�%��d^�T�'ЍQ��,=ӊjռ��M|���ݞB�[ե�9��(͹TF�z��t�9�G� �q3�����\�vx�M�ֲ��,T�О��z�&��aV�^,��Z;��˛���@Q���N�$1Z�*o*u��5f��0������a�6��5s��`����C�8�'�FF��a\��[��]|U&OZ���!����/b("�+,�[�f`퓮�������MQ�.ŴG�#8��(Հ����I��C`[U0��.׌p�c�|	����/-6���,�L��d�"U�ʷ�^L��}�GUNl��+?�ƹ5p�����6��V����}
'��+�27Y,���C�f��K�>��>��>�E�q� E��#]���S+�Z�oC;���RFW�E���>r3���gr5L6�K���8���:�l�-�G�^��~C�@�������˺��Key�����A������_�k�#U֝���P�񎐊=�Ć/ژ�es~���칸~KAY��arfs�\���V &����jzm�󸿈)�0eZ7�/Ƿ��Ͼ��C�����'=i�/�=���\ �Ө_MG��nnt���HGxC�X���:vQ�БXͺ��#y�|�I;D�^̿(E�N���aam��hޣ�[�[X�ۜT��y \�i	a& 2_������$�ݡ������̀,�
6�9X*b���������W���TN{�_�)�!،�����5#���J�L4Eq9bY�sU�rz"Ϣ�Vў��Q4�R�M�.�õ���pu�Tk:+�P�Q�K�L��V�C���!pr?`!���wv,%X���*=4�� �<��X�Q�榄��	�8\-C�1�Ӡ��_v�����!��.�̉!J�5-�������9p�����/T�st0_	!��$�/�Vk�@&V|g}	r�Pd�ф���Ȑ��e��k�WZ��~m��\��w[+������um���@3z�`��B�8�y<�K����D�R�U����&n�g{�G�44N>֘o �*=���1w!��K�s4&����8��ko"^����J4�Ȭ@%A�RS%��@N�[,탟��������f#@ x�����s��>�D�^[�'Q$[.�y=�6�a��]�>��д���Fe%B�GQ�:�zG�>�̙(�KJIW��6�o5�'q��������&G������ᬬ�sJIA~ȣ��E ��D=?�E1�@�ȵ��h��b�HPpƮ^:֨+��_e �Ã��R]�FZ�}C�C��_�$�:j+T�����"�2O��t�/��6��7JPzɉO�:ɧx�./���H|I�=]7��YZ��vh�C�K�0qP�P����j��Y�w�Tݝ���v����������X��E�r�*]q�9��|AM߈,ݼ��FL��j��)�nے/��_Q0�)��Dc`zQa^�f����Y�2<�O[��;g	d闳���ݡ�a`LoB]=�۴��1��q:��E����D#O��]���n(�o��� n˰hN%:a������c��甭�5UO�Sj�n�jŷ��G���0,��ڴ=lc��~�e<O���	���tI|`����t�SVGIa��Σ�����6I�32�NΘ�10֒A�6�ɕ�`e��^Ѓ�X��5>���g���P���:82R��(V�D?��[v��8&K�ȣ8�.�f�kxŌfQ�R�֍�zu��1mC�<���5�x!X(��=��调p˶R�3�L���Y��~�Z]7�͓�&�Tor*������� ��p$+�pnV��)Z�R��ګ6�E҅b*��88p���o;����.���?<d�_F����$Q�`�@ȞA�9g�kA����^S)t���∴�v�@T���4RVN��4W�����g%�ԯ�}�.o�
|���������h���"E�A���`4�z�v�8q��(��;+M,��[�R[�ZEј� ����b�}��BD�X�c����d�IMxZ30��J�n�D ��Cl���	n6Zg��x�{��$c���Qt�[j;\��A��Ģ��e�4�!�dH�
@H���X*'�����^٥i�-��ߺPD�x�"'N�bsK�Մ7��&���5)���W�?B�$&�DB&˽ `^�CO�&����Ԧb�}�P#�Izo6S��Թ�m?�'97�6LG�CE����ϧR;�zT�f�2�A�:5�m|۫��ҭo+������,?�mC!��w��夓�,��|w+=i��ZclL�V*	����lD�X+�t�!/���:��
]��+�Q<'�&���IpP�m����/^긞l��O����H|jY����ᠭZ�K�i�ig�k?:���#5@��N���m	$�|μ�j�fn�R|� �%�3��f;�x�mDœ[��
X�L�r��.��R����N���&@�R$%\Y��)Җ���^��H�=�NWL����{�J/���` �FC�o��]�a�U��ާ':K��uۙ�b+ �h�����o%	-LjL�ůuED�d��_�X
���{��CK�k�I��C��Ŏ{8
V�5ʉk]Y;��Y��Q��d���\hT`�!���a�G)�8��qT,�A���������kWY�]�&�ʃR��B-L�z,�%��۳��\��^B��������_%R�IZ�{Z��/�9 �<�Y�jq��L9��w��>6զ�0}H[��*���M��:s-�E3妒��f��q#��ة���I���049$�A�7U��~����������!+�I8�G�&��|�zc�
��V�[��b4��W���ֳ/���L����\G����;x�Q
��z+5d�AKþM�]���"	xt��5Ȍ1Q �X&4e�j�����Pҏ7>�љl&�|���_��h��`S�"w^�M
�a|x#����iV%ɰ������YPP�zh�<=�'k�n�ĸ�w�&s���(v���B�_�@�|�:���)�.�;��0Y7c<N
s%�=u�#�_�<����v$��R���͛}�Xd���^��SC]�i���8a���®~�S6S�+������O��N���P�m�{�I4���cT��6)� �5?El7�;����ϝ*<|e��	q�A���&l�m(�ؕ���7L'}f\҃2��MEēe�+�c�Ӈ<��?%�㿢�&�;�Q߅�%g]&
�WC\V�$�*�œ+��� B��~���ǽo�����q"D�K��x,�B�q��+�]N+�����1=a4L���JY���l?�C��+;r)>�KZ�.Z�K��ueDn�b��5��6;���n}��)��z�k�l&w��*Y���6��hi\���]���wH�*��j�k�<CE�Xį]B������\}���՝I²3��QᑷW4���b�79ꃐ��1�)�è��e׹��WRM[-��� �����8b��3Lk()�$�3�X=���zw@�5{D���Zu �����@��a�ͽnw�)3���ܳ�"{�`�
uaXKl�PH��l���yG�