// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QthRBZarjBWESkMuov17jlm0BqZypTkNe7EIKxWdBdJrUg+tvMg8ohOhkQ/+X/pgvb3WoYSG2hae
4/YPT1ezoyFgZcuVX/tL8NTOJUO7TB4aol3m24BOgVGIS9D4CVAEYGVNsrX0h4YWRHoppFs3/ILz
RghQfD4hbDQONndJlfXJCJMAadJjiE+2B9RwRRpFvRi1eCL/YcMmNQmvdblvF43bCeGtXhZZ6OBU
S/s8Bk47U+H1CJfKwduK55MXiI6oscUQcyJVmenblVNDcaKrdetU5e8Q3d/fnb0dhc53Oaceu7OV
ex9nHQ2lCRTL1fNDuNVPoyF9ovc/9sfx2+NOHw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
3Du2aPABoOGU3fRpOK13hg7aYg7gbS93yn4hwC8Amoz3BRMAye6RyjHd4icsmaUcrlX/XBFX7rb1
iJhhEpPAIXpdDaLfCj4VR5Z5DQ/9A7dSEuyLryXPRWt2wjaYFV6/JmdYhhfeQ2IHBXnbF/pxfBVu
e/g6XDSrFzJJ8Cbm7DPHX9/C6LIAbPkKHGh4shx3M5u5kh8C8AQ7T7Wpjzf/YiT46H7xS1zXvAnI
zDr3Mp8t+9nThaBHRDNDy2A/zKEfBh6iA+OplED6wbRrtNJWm2f+WpgOlz29jqkHhF48W80TRmIm
JrDhdyGNPdhzzS/nkFVF2CSI03jS/OUDSNmK1OWSoXxcqBQCQzDWQF0zo+DFVazW49txnLgtsutX
jjGLqIkn9ZQEVEC/zi4x6osMLCVZsoh2Y744vAF2rqAspMZY0GVsuJD0vdmZrBJsehI3FP9mcgDu
SP72FJHXj+J8hsUH3gRzP6z1FBFzk3eqjrNWrM4L05Gwy0h9udeLEZqP3mmnomGOFh6Ux6urm8Cv
Vt/ZOrwUrbQ4CEYoGQSbKo6sBII1RR8skFC2nCzyNSuZsgSgMGIIFc2eD1w1hQkpQxDhbgxtYO9N
NXcOzw2jQMoBptfudpBjMO/w+m7E3d+hdhKhZwUfID0NdRtkOOuVxx4pkhwHdYeVJqxBHTxTyTw1
he6WlZyixf2Y+f7tKt7przhLi9BKnphgddcPnzH9xa+41wPjSAR4HBqbdeJMqqgsghbo4Bo7lTAO
Y9vNoAp13e5kUzClXS6KcV2zOooasp+W1CYUyif3AYfWG1+k7vg73rVe39QT2nRFWj1XDhG6VXMH
YC9ada2S69JhkKA+dyESdvkzSf2ldnUgTOC8OVp4T1cJKCXW3kE2y5ig8HKsbQMyZZ73Ni5/ZCuw
0tvalnRgl4PXbTjbn9N98OsMuhQBEFFkGPXHW/Ii9/LGPtQ1OoPtRhS5+docEMXHP5RB1+UoumlV
b+Bnd/njK8OD/EbFfJqIRJcO5GWryEAcqPSBd36RIstyx1HXx6vACRs7hz1W+a1irbiPQOJaNwn6
oULmhP4eqcVob8nS07m9K/vHQAoqLYCyXdm7+xodOtn+176uFB9McMP8SXdCRh1cByYT6tj2efxK
7STWkbKx82qkJCa7fHtFKc32b32CN33b4Y0/BG7Q2Gca1/zTw28LMGjX+8tkcWk2xvaOuXnzeaZ2
Ofhob64/F8uMavsZEf7ZkyDlgySgSWy2c1q8bb9cULqGzgZb1tv9UjpiMuiopBwnuZjpKsbY+OKa
Lgr5NLTsNjXhOWhMnCjizpo7ZLWnlqrTEUzt5CReKPsqrYebqs9YrjaWm0DAYXAzKcNxIHPSG+Wi
zOt2m3Dm7W+c55WR3SIZ3UqLiDAgTNEggfWj08b3CxmGYrgusexsvMFB5FF+cghqg2ElV6HgufQ5
d1sDyv0VQgzlBQ5D/RTZLoRjFoQ/ptKSrH0X81EmJqCZ6lyyxekT0LZfmkS8GDGnY3b2RN08peDS
lYp+cBrUAzAGRkUwicVuJd/GPxbOuTYz9FJPeq6O+7Bs9aOokDwMYjMzk1dQACBsKi4aMBD+n0O9
4ArMPewoOW48Eel5vyz6mEXmXSxFeENW1s4uS3cO9HNjOIj7NPjaLkNYdH8AXL6DA1zKU3nSGNdD
UiqwFwTbkKLIIbrcYMuA+gv4eUmxd9qiMcT8wQL4PsseymXDYr3ZeKADfxnWJLAhaPPA1x8B1mkM
G/Ov1hwOMblOWJcThc1S0wVC3c2WUnc57FkI0wRCIdRkeXKM9KOmDZ9rrX2hab3Nyx9UR3vGjYJc
AOKvccQfDJGinvJzTvKESUuMEqwMv8meDwrvQrFgJSmzh+w0I4wf2DDMt6REQT/L6G1raMTGUIaa
q53kbHvX58bLZ262+HA6ENIA/cKCI1cdp2ESnvpz/Ypt5Nk+kn7Nz75VA4cB5AtX8JUCBTOL02iz
wnIwP8t2PTHZ/KN8XA2OtMzeaiobD1bHYmjL1tnp7jg8rEtS6lermXJ8XSWZ0MCdnhkUiSOy1l5c
UCY+KkSfZz0icJqGgAplkUpcTxaLNWrOlzlACycdqyw8Q/iPB2GKkAvnClYOU9hgqKZ+epsFy5RL
4FW91fMt+46GFgxRQS0rZBhjdRsCjr3UF5Zi2wtlNi211eKFEFAdPbwH897UYiKk40xJWVu3aWaP
kjx9N56V5qH+1BB6lHLg0Abm/Xc5v9BSEp92UoDW/pSAA++hTyqz0PespT9lSMxq0Rji2OnhGQzr
SWeFToIPPxtm1hjKw/snpYRO6ej1Hd6cPsZwxnqq0dodGaWo6dj/WxScUK5uG4YLWA1QlpW0qOFg
GDErCHO59pXzjQHkbVU4VvUj0Q5KxnQ+4waMrblJMgTyuTyr/s8rNgfcHV0h7/Jl+I2u913tZ1cM
juxiXqQa4e+wkB9ZfgACzdipjnZ3Tb4b3GhgXm9p9SO1shitSi3DNtisKVjTdnZiCNb2dPVbCIxV
sWNpOK2fAFt1QcOiO1Lf7y22znC2xJXV189KKOF6oNiAIQxZ+cGfbiQCx+JMbsUv9Me+0O/K8TzW
F0L/XuBzFEYDi7OlXORlVz2USOrXIgKNH3vZGaZq5CyNTlEdXIvff9MA0oy7IyIttMK9TL7aKrN9
U4NtMkJozChI2QnCd0AKmkBa4wkb9BEWKiqtQFrriHJMW2QMhNW+sNwWHXcizjeSeqxQIJy0baZ2
ryjSE4SliSaV3Xafh1lLTtNt7YYM3IKOKpArcZEsvX2V1qebiBiDpaPL7jXB5AfjyFMZtiqUhmF2
O51wkAkI5gf8N8j81pcPrZXKA1KP8JjLbPdly1Lrhhp5C34DlxN38LaO9xYWwlCwzJMKiYJ9nfaG
YJqs/RSAmCZpgeMHHssLoLYO+rE2FYPwv2wZ0ki5A3Ca5sCcETkOcunbXUPLm9frRkyLeFwyOPnf
76WL/Z5jAZ9A+WQaII/IapxPPdSHzg5ULBZpy0ob26qiXgWXeqg7fc/nkxUqhTo9RQA0GSbhWPSa
+CMs9SkP+qIcTJHMArXgDeNlHpvxOtVgYSVBSSUro/HIxM7tQ4fT9Pnyyw2y3itTfgPcod+BLpQR
HYCv+fhPTsO+F6DLhkeIi6KMWP8rTsvcrOMYaoL0u4qzWdI6s2J+fiPDd4gul9ss8EtGkIOAVs1R
ewkXoC77J5PC7FfMUqVZs/au8X5Mm1KwTZz5Ga21xYR74WPVYu0UvzVwsVXip6d7PkJNY067qZrr
PKuroJ2Owq6iChU0i5osL1cQSq7UkxyRYU3VctmoyY+f7sV1BKp95omvBrdawQG5DMTyq90coSJA
s+stjO3JMP0Zla9puWQUy+tcY/+vIexIQ3Ap8r1FE4Dy6CC/coEfw56z+PEw+4JQAPruXhLt0hJ/
mdLZpJ/J+ENmCyUgqUFYvstL5u9tArX+kOXGzCrTEhMBDI7Vkz7/s94DbSdEDhMOzcaCLFVZzBv7
dQwwHJjnqtUTQjhz3Gvf+GP/DyRGpKO/VrqUUBUY+2kfBMziEDScOy1YVda9bh493nMTexoFxWDv
4ZJB5wEEAd8iYLKUQt4IUt/G/tNV8iwF51RlsFj5mIrttZg54t2OReu6M7q2RASpce3fUcznRuMn
M41ZgzUwajM7t4cNH13tKlqsunEPCR3+kSY9JTBZKxw2q/dY23xudwttb7X85Dx7BDJaMdLMUsEs
YwyxCYZU9I3qcYlxBuafDfEkOUK7uEBsrDrAQN1ZyLo7vybW0apBHTX7GygxyWw2unt/ntdplVuW
EYbM6qcNgEjuZIa9yZE5MdPL7i/ekL5Ln4r03RLeD7LXnXBebpRLkgoMnA0QyC7tQj+pUb1GOUVw
/uccBeVNG81JUm+JpdyNRlbINzx/wBrsS8wvuo6QgEgUHivA8XIgB/mOFJmIiy8aAsIMsAIf3JhK
v5we1FxgdU845cP2UX8FYSBD7Y4cSDYiWMoj0x9Bx6HJ9kqfi1OIEIBhOqPUM18DxP8FOXb/SEgu
68G7Fyqn67MPKLpooEMmLSwkVpqsYZdk6vQFDxjsNhleD1KaOfwLtv7l8Z/c/uCPAfUJ9KJ690YG
7PdLlkxCsF7I3txRk7SGmAAugM3RUafQKgRbWX+IjZ0Yqv+D3LwJFW/cj88UfiKY84MSk6QagQqa
Fko82HawzPi4vt/JHWKXj9WupTO4KBAyrNqyak5bQ76lLAQEIrR7LyLx+DLMidecY955pY0ZGQKN
01AdI5d3BesxQ1lexwHihznf0zB2xkVyCSO4ElHpf89kV6bFMLE3mim4ls0dfp+cvFwPft+IgJcF
ag3DOkb/Duj+svGzDueY6d6EUmOavJl8SgpjXs5Ycun39cY/VjvCI+eTQpGGQBdzKqEouoR9MHUR
kU2WdT6dQA+QNXrweEStzJTcUlpGc6eOkp391AuFAIHH5QUy9UsYBRa1AIL+D/V7Y1nboXuAFXb1
FQwpf+1tRBJrbnJZCDtfopp/Arl4R75uAhf8OFWA2mobog2AtZwpoiWqlhFdSyoRxxgGgC/bV4Lw
Yc7CJAkx+0CeR46nsN9jr7QesDpugIjfXAe4eodhwYhacrO67o94NRmcMCPi38jfdwIACD+Z5hQC
r8JjQr6MOXsT3rKfzrWfs/3NnoI5Asza6867LiclOJ760oKrZ4CE5568ljJxVs6Eh1GHLZguQf8B
7JXDfPaMCB3SSPnVIQkiRzvkoXtge+cGmXiYoXkEj7MAc+fHOd8rhOTF+By/WiQU6SGfsZuSDuAY
Mi9N9+1U9qFTlTVh3RRMtA6GA2HCJw1ef0kcmLoq9K/pTka0HVRbYtQSAXbG3B2C/yL/6Ozzxa1K
XXp1U91fVTsm1Ytzsbvv5n8Bwn3SNyxg7TPYX3yT47P+hYnzh3pW0lmh/+2Eqm5wbHnVSXVDrUKm
D6ZkHenhCthBp8nUh3jeoBVDsEuCJ45BQZSP0toyzmx6OQiC2WIB11v7332RhgA+1857ESqvI9Ba
/kP/5NXH/kPwziHzq1bph/jWGJVa94WtC7eBz4deZpFEs4nKZNQTROTfeOw1oebsnXkH7ufG6xjY
sYzF2q8pRJiHI86+hj5KG7yQwQhMd3Nsp6OZYsUfXId6vEsdF1Mc1LzbmMgPGjJ8XNKXrgPGyHeH
j5xXdNgaDO8pUHTGD2ITOnFJFY0oZNOpxXMNpzKH9Hn/Dq+BqMUIJKtfz4wKX661z2/YzqUSl/FN
Oe8WXsVd4iBdaI7ThIDo3Pm+aLKnf04B9zHPlghITron8xgEkmOxuIy6pa4KLh3O7gBbf5zzqKen
Q+q6m7O2Kwjx9A48EASsqhSRahAOb5hD9KfYgGOlz7x/wXFDBsk15BGr4LTiB+NR9pn4/dBE6d+2
PXnzLCS/oQc6CA73tppJ6KY8YDBToGjRpkJeh/lMj+R6KOS1Ohb1KbdDqt8rbdsYRtbHgOWDrt2g
I+eZ/XlooGMe8a3qSxfuGslnHpr/1iER2ZCLwt7owSi1wkTttl/8x4qkXAsbFEOALFHfq81pfpxj
HW+cuXV4Pe12PCuk+gRutEi6zEslu9x8R34OJmulzQh+eEdEMK2c8IX6s9D2SIsKhsQqRHjb7TeT
oUSB4w05zj1V1EayIij5BWAtUoyHYxhYBqHOZtWDutmsEJolspFf5TdbDcUdGbeA23p8RqrcRU2Y
wFLzdmPnd37NiUWpv2zmhb5+VhYFPeBigng0AFuBKd2G6XDbGJYuly9lzP5J3dYfa5A0AMlqduOc
TCUBg9SXBRy3iBx22txMrS67mAdkmh6WkrNvLHl5ozfvwQNTB+aubLaZPe6I3yG9Gy7g+shpa0C/
IRThObuYIPwg0bc0LWyup3yo/6rBgOt4V3/6SLbTNdUltl3y8MrJOIZyRvrkWr2EZIFeUXbR2ALF
msFDX3cMY48EFaNhU4UC6Ni0xnIE6+UdCKTXarRSXUsuh4nYcEFmyxWLtRPVs99xN+YBNh/cEE4N
H9rzy2MNnOj1dl4fLlLF4MItCD5s+cXrbxIv9lSXQJOi5HamX17Vq4gDPKFNLk1c+St1S03ajGLp
chhLkVjGgCCldFIMXTZ6bA6fYHj9y8LmqZmw7Ywsb1nbWRzwk4DmnOVSRDjj61LXzfKFXhLVb2y8
BmFMs2OohplBwVwBLTo7WL9/GXcQ+31IEpQD8bqN7/1NdheiaT15EHR1nyvkrPQOhjC3y9rRXCtI
6aMTRqfpYoRU7Lj8ochfc5GGTtUL5htxR7tauBzxPLlX+nUnqNu6/sgP71aJJaCIGbamUvxvozjC
5wt4wgDrpZX3Ebbfq062Q+RJfEEdqM0EBuEuMtvcjt5ZqxX1nZsTuhL4nNT7iAYlgqezB/Nn746q
axo2HRFQ6g9BbOS9nXKKLEoAnJnhIIhfPMUSJxkJu6L897EMPpqPKSyceNQLHBHR5LA7Hz2ia/5T
Jh9MK48xnGxXnCvNPyW/eUw4PSs9FtRahpCZjnJt7F40Gy6Jv+monBHi07C2LfqUBxrOKiDoEGV/
Zea1VcwcUMI9cjxUBNWAPv+beyq1E3fk+Askxfu/zLCQ5kRcf2c6w9EC3NnR7fsI0uS/P6ooaW/z
Ly21KURca9UND6e5hqBdlzCFr+MIzqFrELtdy3XOZX9gLoc/QTACciNl+ELUul7EGlqBzktSgu05
+xh57oAdcaiqykdHBMH4wtN9GVWHSoJI8MzQjom7y/6wvwoYlIW4eLxhB6IF1kiXcFMk9J45URrK
Y9u+AIJyDRfQXSLQGiQiNaMnY+8XW6z5CP0AqZozXGF0wCXaUCxLPepYilMPSYInlYd+sse3LGBx
xNJeQFuxjcEP2uW+YkMjr4jRlG6EjzsXVpIG5f2VyCYT6KbQ/ccKbL+JQXj2aMWZjPjp3Z6JhAaM
RIGA5TRyaOpXHnLrB1ksJJMeydHcgXtxmziRiwEDUafg3ls2BtV3Vqk9DexWC/gZ6B+2v1VU4i0V
ILyAXwap22P2AKs0nTUNeNjtVScATdddLCrtPUX64HsnIO50IR0oR7FmPb8u2GLQpVUVgoCRiomu
bkFdmR9aI+82+BbEsxwAYd1hYYFfJgYzvr7TpWyIGGs/TCfLgleveuhTEtlnVStnopea8WTsZxPU
rj1ZMSC60nUGxEZm36HVaXjidV3SOtfYPEmafL3yzBvQIZChBL++BZea43RmdCbksEDd3hkTRbJX
g5jhDvsoH3yX7UiObRqp1gXoR3qDjgFiDBexqvhVWgMQc0isXTTugXCl7oK+YIRcqmROd5Ut587j
mGG2SYwMOrA4g1BrX+7aVxQUHdcFEWBYP9imlRAlHgBzHJUdBqhQb7bz/lJHdEkot+qAEQrxVAvt
18Pl/yfm9fqoW0bS4IzFRV1ygcdcs+YcRSaeBA7v2U4cXRijOjAKDidelp63D+A/MNtDWxnkdarH
lPdr8rjhYkbtQZPBfWM0XVKIO43cuQg2azB+3m4u7zo0BiBfZFOB5kL1mN2AxXFgM7LOznKD3m61
Mw/7OPjcdgC7XsyMKmkg4XG2sZEcWgFv1Wp1ujDV3tvEKxY926w3Le1Y7wqaGIIiz6omyOh2lyHU
T0hvomj1bA+ik8u5Ap6E3R4OZce8zXaI/CAuOASapMdRbQmi016GSSwfGf1oDHyantgjXbL/dG4n
fKIaJI+Vx2jOraLMcKe2Clbl8coDIRclYkOzrJWREbCbvkUxc2nmFi8AcEdQYhQu4kfWsqSwdF+2
NJ/Jqa2Q3UtxTMQ+5X6FSk1OAbFBn12h5AriwJhWOX/9kjUsiUH2E320TqN8ArnQMY5uxNqy6AEo
MHzmSA3UqhRbECDTWOpef2lOq8lj9S4lQ7Un1qtrEKnHBaneQ9SFsVbHc+eckCvvPkiPQqMw1fb0
QJm0p5SIsNhqsyoVvdyG3Uir827WDVHW1b4qe0xhDUqsQnZ1uj5YncL3MInVeKz8kmUM7TiFFdlk
6nsLXBytp7bUSp2lqyWXAMWkvY0Un0ODE9waaQA8TbCindc732X16hznCLPBaENkCBT2xgrrqVCk
Xc0dMKxhnfRl6heYBiIrhk0dHJ2KUSVXlkq+Em6q8YX/HmQuYNCSBxYzVoOqOsENwJpruHoJo0JN
9xlUEyzSHo6nimMG4BvcbssM3cjMr4YDQhlSqj5nJvZtqqr7zyTiurBsrbkc7XyUeFc0CbQHKVbI
HRvP8eNUnLMynp0cZ0aK/jjDcUTMnSLAxqG3uoUzMnv7UqDULA9DQdijQ+UjSN6ClggXX4eP1WZ/
lrkkrNSrPpMh5dWmKCFQQtWo8VGEPdYkvDk2R4XvxmkpKbwKGJWqd1Z7C+ZX4GJuogQmx8marDiF
4P6ZNGveYzNmY8tC7ikNdzctzmv1OwOqxbdcP5GBUT11874dggmXWSNJUdW0lrfuDvsdTqb1oCY4
ndgyjxTu+V9cY843Mqbtad0XgYinh53bV3wPE8cdPBudktyWvIsj8rYDDN70wP1Kjs+/EDpfv6Ip
q5O6skxbEcnELV/rH+Cxv19tumqOUojDACU8a1RFwIvdrGCpDHM/2UP9cksUcIim2U0BGbd4G1K5
Q7Mfxteh/SQS5LpWkAfMh6i/BkfHuGxZR/kp1QANpDDU1gMTsvBY7G2fLj2Y96mJZFpcIOIHrBfD
ic3Eh0VniZY/igiiyKqgsDfwXWj5FNdsmmf0dkiww01j6E6Sj5wk1iYI6Kzr6MZ+h60K3atVd/f1
QEZBYdnErWfxwdISf1giLAoI21/M6PMgPQ3xXabxV+AUxwLNAD6rxsprG+nVZ5SV/9zlM0n85N6G
EELJZ2q2u1bAkcGDGcZo2c2S0OCfNMHbvEJwZm8p0+F+aQ4R7cg/BfCdYtwq4JdSru5hPm1njiWc
lTt17H65BnrPLwoz6qJOB8j06G8zUpYnXDlQZdU14I0+D2HST5O86JqLP2OXeeVybvMDpK53Zheu
19eWvj/zLKsbwrKytstLFvniaeDdYcuiYZfi6IvYlZqdBpzG7xuuIOv2trMC02xGBp8TFq6FbOje
tkbO4YDWAKJtoXFmDUWWbVdEtpye5jP6i+XL7zopYGRASSCGTx5qw4b15Q+jU2TM0UUsJBU0mEVg
MFLCOKFjXAymmAP3OmUfS0X4BL0CA4mNmtgHxDKHJnK71cOqp2arLyc3IUG1Z8gqtMX5XaQ1S+rR
c8TUOYwV8GYYz1UuZMoPC1yh8npUyVuCZXKPZyRi9ya1ia28+bh/TSFqVguuPb1JFnnJ/ZPlhAck
zoHzvNAWQZXMivB9+qKn61jYpAMy1Bd70BzIJIlSPJCirx7P/tHWwnJnuB5bdnVCwUhxVNzRykgM
KqRmxvX8tcqMHKr/JZkJd3FhYbDjnEweqGIdFW+0OMB4FR2BcHue7GLFiLFshCzptbChGLNcRuBm
buWnvFsqjkimY0suaqO4eUN7Q5n7at3gE+u34iQP+B4kSVgOxX/LF79R1HwKlTCPI6eWu5k6BTZm
iBByjI3VJYLOmTGrVYNYQbRjlebG9XQhzMlvfj62JGQz1Z5Gge6db5FRxhEdyJjazvS/ZEUcb8uK
HjfHByMBsowV1YLUcPOkfGePwzvaAz3BhJceE7Yy+ZaKaW9NwVrIsErNtTsr+xS7BUkKW1qytC9a
EKIah/xITXPMV4ZfvxAFujOnK+Vn4i1F7Z0cYrQihABck15qM4EVDdVIh+XaxyGM5Lf0xpszeRq4
SXJ3vsWf+M16XrPkPpLoJtf6JD9BtwHhEo8UD5PWjrG4JcxdgDuoCRPQBGTuTZG9cqDWnjSaAKCi
j/389fRgqVVqVMz1+rBGmsWiRTkskFIP8T2fdXf8OYMzvaVOYyJnqpybniRco1EScpEM7BoySeRB
UdzBATXdk5PTMV+8T5NiaaxzrPGH4l7BI8LIep/tRjDNWe6PHf0lpHDRMPGWiujmbWfnxYD71a9j
6zSzB/5GBuK+vpgyXLzm1ZqJ+WMyqgUbnczzRpOQlhYECR+q3bP2E3zqdNqPOp7pgnODpCgJ6Nx4
FkcRqK3fpud6z2I6gN8Pg04tlJSLhv+KQSmaPCMu2jguAsMpeaC4o6Nys17AivOYlpnCAir9CCxQ
HbeVwuJAnU8PRFv9AarlHDCdDnjlRqMrlVjL7PO8bj7xdG4K/VElYvPBeIY+5ySQKt4YZ5fVHatY
veexKK88i1P0AXxFe9YFf8HcgKwPU3jd3nB5A3WHt651mCcr0NJG03yzlPRNte+EloDCO07gLWMh
GG1EpAUkbR6NU/TcFWTO6t2fQzwUMD3PowAJDU12hLYZKoP6vNCLeRd9RMGueaUDkPqKLOzSLgmn
TnQcGYZf+Q+OJOakPO5gHqAMGIxjBuDlNe3TeKRm78YznVbzjKOZ4SJV3E7yGA6wSzvY0tbnOt+p
NWwEzYa/a696xaNdiAPCapiW9tMYsN68f2TE3Ru2bPeHAzPAdIwv4gINBWpp55bqwko6MGVi1YQh
Sc48eZWKt3Ioz2VXYcMzpXwHiLdH+yEjeCk2lPfkSfMc/3Ylv4gwpXZJ8n8hXNzuzzLMorftLglE
3cI2ISLeJ0MvOKwWozV0LAu9YyqhDt5RV29rUjL9NkaMOYC/RNBoM//jnsI0UjiSAcG69F7lopSi
zCsaFpdVdiyaR2MjX6OCiUqs9ToMo88VJW7PZ8pQVAljGo1T49HQP1siRLQwcR6y58fd/Olkc2kq
9+yTstqeHx5Wi7P3dSfdFlQB3wS5tCp78zV9tCMwpVwRRRIrsosNrpQPFXArxD5E6tx+K9NOiatB
WGtb54Zrsc5DSgHAeth2rGJU75Ubz16BpI6L0s+KULv3sW5+rPtPjEq7wH4X1aABWSQhoyx5NqyT
00wQmVWeqoKgCZfgccEjOrTvpza6Dx14vdaUeQ21Rh62LLGGvFLjOszWD1+j6bd/P4VpfSBfUfFQ
kVOP4dw9XIjcKNbo3VWs9M8cLm3lwxtPhEy0aD6eSpCUe7tVbAlOUMQOKHlnJ+wOlT5hY8v3FGTm
m46aFSOpZpZn0TzNvr+Ov+FKXN5TkKGtRrQxl3I106UrIm2eE+nGF24vYS7H6NhJFC5Z/918Dju4
Wv9+JSH9uQXNwN8hkgYo1m/UkzMmDBW2Of/buOt2766sICl5jMOKKd+XT5uStXcCx1NrJ6BJA9B8
e9sx4ExKM6wU7sOGFBhhEGpG3f1akOucwPUlz2hl913c+5Ks4wj0/L0XM3J5rdZ/8ZnNZiIEr2Lk
QSvjB4xANrPgY6OXVrzwGWPBOPkbL8Tj75bchCAozJp6pILw4GxruGqyRCZEAXEFj42Godpoc78m
+klWtH2+X7ax/evIEMrN43jx5MOPn2P1hm+Rx2eb3B0WmbMPE2bHXCN3Adz/gITvjLmNo8qJ5U9n
PdwV8LWNL+ZaGLZL9BbBQE6vU6vqxt/fu+Z33MirNcEBXG0TsK3DzBDqlo7ufMJiVG0+EGBlqOfW
Su+FKI37RUJ7b7TfVJdmD7PfxMezWMrSrb2RD81L0m5RSKdZYsYxXm4EIU4504LECYEw17DpLF+M
7PtKN1OLu4hGVyRYSTMnQ4265Vs5J2S27ePPDHPul6btwNQLi+3RwyO9CcnGTKmLVEMwPwz6mPHy
bY9sRxKLURoySjrVO6VaeaF3XCDtXW4y/5iNY5wiatn7WA0Gyjbt/r4ULtIiWSrOjgvSIr9WZSdj
4/GLcjhfHLe57eZwut7YX++wqiXorfEkSLuqqi92bYp7WcUfEThj1uWxf0yc61j8fbdfGGLgOeWO
GPvJH7leoFwKhW/2fYrSHuo+oxqJVu0CdQfjDCM2bpYX85bbljIFq43pdcTjhKAwD4YE06WEHdfT
o1Jx8sZXJJFJNehMnihk9bqhxNzPUDFV6F/cSTfVJf/YKqXzM9fzIS6FLUIi5/09PNEUsVu06TFo
/5iWQxQdLvSx2SQiLcJIBYmpRTBV6maYaSOU2xQ5m60jLXmib6uqnC4LRRMhVH/YHo1Zw7d08vwe
GYqUG9UnpStA/g/Uc3sA+yerZX2N8U8hYD8EfcnnXmPtTmeoigV7tKrrjjz4ZRDXKnhbvPGepBQb
b5WQXpCTXb8Gd6rgbb9tghV1jpX6FUQori1u9YdhjTYTlxIIVKnYUk+mxBHY0om6gK8KYoBeWVhU
U8LnAQuWdyJN4G4kpZsfTfsSLnOfXtHua2ZHqezKkWhD4ZSVOjAY+Gid8ohiTE3Bn3aw4unDxoCA
xtOMMMUHR9adUrXo/55v/wKmmtgjHZayTmsRQatoSi+m5NwwNXJtptabVhBDVnP0+sVIOIM9D/2f
qNx4BO8PKJM8RlAh1ZKZveZ5oJzdceEM5EbvZEzVLbZFYV9DjR/qHeChMSMmrS6jVchBXR9du25s
f/2a/ZdvvBuiuOkEnJf7QXuyvyApLf/21nbkfngFiHuYbVFJ8jJ//COiA4v3RcbU4Tq1krpRhZgu
h2SmjXriwEvgjxYnDhfl/Mj+EX4EXORJLhkE5IDEir9fqS20thyBBY/mFWLD5SN68hiSt65TM5kP
8sXjKKJpO+jvN3xSYDC2u4i0Fof0UMQEfHnvI85q8XPCWk5HhIRf+Hho+YQ8NSGurqqGtYarCqEH
5kt/m04Oa59/6cuDYU1O2jr7ZyYDEEsSXgnGRcytXR69wz7WMCBvpE/YX8ZcGsh3FOTyJ7Q0drEX
ThNHVLDobK/H0HUetXYtsHqv+XPbHGgyDXBab63Q3QRA3E7OB6FKv9ZczVHh0+8Hns/P+a3fzpe0
23eFlu1gtlco9k/HUBpGfG13evBPPIPljvXQDMOyamm4T5aWFeG+wkiVwLcgWqPDgab5yxEXFFK1
IfV+Yq4T70FAseUOtqP9Dm3G7TI5+a37ngF/7YHSCapNGyzxU77ZbpdZFY1wqQN2YNtH/tNYBwBZ
iHPddWKEV0yvt0UUxi8RniwuAQRvb8OJLV5s4f590uzGEaHQMX0+6ipIDmo40/CTfMmu1fmYqG67
dQa+b/waI+GCpZob9guDtvuMwLDezbwxiELu9jVc1YVM9Xvnx9D2UvtuwYI2t7wK8VPt/pgp/zYZ
nKmx5QJ7CzwPH96cd0kiquI3TP3p2Qv9h4EIU2CuGv2nMlOvXP29hdofvb/IZXuRTyDApyx/SJQa
MNGX9E41RCgajirGWAjnQqL+sZtm80Xqt3513fzanMF57bWf9Q/QeK6FAr+O+tB50/DNJRNBJIy8
+O//kxM2zVwsqOKywrmJi5VXq354hz0rfV33OkoO5sGqCJjJsbkDtsnL6aXypjiXw+kIImtN+jms
0H/woW0OMZFSz9ksNQwi1nMieIrzwBfArTk55Wh6hPiPzDbJ7URi/sgDxhiWC2bjqgCTkmJAmiRD
5/OoH++LnXGBxRxcsGyWh9sHC07TYZtclZJPq0Zsh4AYGJdZIeB1Nt1lGnHw97b8xshncw4hljVZ
COMn9EpUOy00yH5U+c/1HqaVs4J7FHasfbvddH65ig8nw0BGwdL7Nog01t6TplIebPxpv77emycf
QmqxkNCVFBpmWhrEUutymGchwvxRZs0Ka43wxY1OHjIyfQWJmAkL7zqok8AT4oXMvZHoDwhLkLzy
e5mhGYWypoU7HQJkVJqZt+zvgy6LjaSfWsujURjBiB8fvw6/PgmtGGdCmupIie7qmuKCTpmY+gwI
k6eZfrIbXlNFKQ3+CvNJvfNEYkAHI4PCMii1kz0qoQyiUJpVIhY/xXEIe9iabgZgj2cLym0g/eUl
qAlQLXALWBn5AM0ASLFq3wFwc4yxe7nItoDpXycb9dkcRXBKgRBJzyWnU/TDssqxJkccTX7MJuj4
2Yw58ge4nkadot+0Xd43vuX41qUIA3AT1fFwSBmJSM/ebUdmPh2kWBMUvsTqinWIOtZ6TcZ9VWWi
6Is7c8Q2ZWRbegopXwpbYF2Hoq44mZr8/HOFXvPMhw9/ZPz/d/4J2v6g9GdDUJpgd7Ddbj6dXHDA
4o8Y01i43AUXpC3ez+UYpTpbfrfiCgsKOY0mrvVGNQnlM6toQXob23wxXL8Lw+W7XFAPHFn9Z7JT
ciSF322s0+/4ojyUQelezh7UeWnYh6Va8HMqXzxzTGKxUlpj75iO2+yvGjufPLmf3Gl5p9Qnmmxn
B4gLBZuXlk3U3BT7T3zrFztfQzJjm8ywDFl7TUgqGX3OlpOlm7IptOh400eQlDH06/pzEEDAF25H
UbPdSj2jqqqNjF4CYXSSNqmitBNj7E+c++ZxkIk3fr+UEhC64w28+FwbCSMIo6csuz4Ufg9kdi+k
TdrlD/UUqrmoROOIFXbsNAGkebiefqLSPxJNqt2q/HupV0G+DdDHXb2CI60n0to7o8xnNYfg/HVh
ZoueX0dnHLPFoVcVhtmay/hWX8wJDKqCaY79ryxymk0T8LzENxHaSiNYJUi1sF4oAnsjhTb28gS2
b57/luufgG2/mbhXF9FaBCM5kl+Vi84YeGWAoG5LI6DdGb1kMgKGJ9eUMmWJBS6/h0tkQ/3K2kXm
Nn5o6ZtAncjq72VxXT3+e2Mqe8WIYcKabUtxpX3lCkmydv77gOIva5usWrYq4Nbl8ngzx1Pu+jdG
fF/CEKsbGnm0I8/Ilt+RBd5SyQpErR5xAegUPJ3eIu80Irdn9znmUYWcZNQWxfO7R6p1fF4nylab
R/Y2daP65yy0WuSLh3HrIEUL+6bJ3oeDv/f40vHbNXgkKAqUy+4Ap/0saC8il0GPwzAG5yAHujXs
prrel+Pm807Bp6Y+m88WD49F16cgASXz7ePqSzGOH5mrTec9kz16St2LbTKh4PPzfDlFj7JXxaCe
q64BVWw=
`pragma protect end_protected
