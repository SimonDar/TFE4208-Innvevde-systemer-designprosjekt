-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WdvqgSX5MlPKcxNA9YBojMM8N25ODNJZ+bP3RCARVR+A0My1hTMk9S2NmhApSL0xERL3fnLV/7le
YjpuHLOxN3P21qBMRGz3lLuER5jIR+5+KadIhfIpJi7gwQQr32KLlntWlWevy0DhpkRnqr+rv6fI
IAS5ZYBuXlU9WSBBBXnj9r8z4HdAgTMXW4ySznoZZa/pIrFtXGgTmD9wfYgC0+OoFouZITXgMpUK
ze/euef0IbWtR2J+Mz2vY4H5yERZP4XOPHAsvScnbJbtGRyLFEdZxQKn9qb73//trps6Iy5qiqVT
nNg8AIU1Mh0sEZPo0rO1wpTHIDAKkcal/TBvFw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
pFZXdIXCCA5gPOstjN2Zae2M//WrMy10eRAnZ2bXR9WTNKjZjDko3TQYUb0WkURfwVOTPknTXQ2a
IYsy3CREl7d9m2MbpbJxk/xfzJ8IiQG0h32RoHoyzP2ot53cfcsK3fdUEqSpclexvW9aKZptKHxp
JdOBVrwaeeRPGboiPko+7Uph/qTuQLu9ZFsBBiPCNaexVdawOODo7n856X2qIIujG+kmcNSF4bIH
ptaWLeDyJ/38LO2nS9hmUHK7wM7l8JmRRGi/0aWxDx1RRWXFaEhi3qAZ6Uy/izbn14b44uUTeUAq
/SzTQ2dj3G7VqlxbuOYnk3O41OeKenJbPARQaK0nrxw9poMXGrFEKXf2VqkIYwxv+yTAGTofbmz4
k4zIsovsrU7qZu/Qei2jj0XjaN5HYwESKC3G463w8n2y/CECVSdwl9OAMA4rJzfYplDyTKEXJz2k
cYPRe5DzOdBaJa5j42JYPSOqu2ax5llhHQfj3/9WcLW4RX6XTZeRKFarzUEwAOmLfl9G6NshOWjx
MX0kmHWinoH7z79LSB5wMU3YB2SAuhZ1Ar5O+yhgTdp/pHws2hxIOBpKlQyFphlDRwWK6q80w9BR
mqxU9V5l/R4avpOUbR8Kn7WTSkXNofs0NXCyikyqoSNWUH3b3HnsrmtLH98vPjjyEPkokihuIO5U
f04iQTY3uZ/p5sjDX8bdig0zMcXrve/FZLXmX7lEvksecKA7bmMd7bgzfb0ic3CwkiB3cryjxnzN
w9jMSXeaIIkOHcBn/6qNpKvKCnh2ON3nH9wr7RtMiC28MCXTFz9HU6So46IFao8M6Rs/6qsqpnH/
BkWAPvK6l8PrKcmb9qNFrNzcyp9mwMBU28Y4e+72U5BZn6+FT6eTsW/Jpy+Oo2v8YkYbymP5LdfR
TaA44GDbIgm99V+ivWOCIjXHCLVL3S0VKf+9Xmj8L8dIGrhY1uEnNnpu7n71BD8nN0mOUfJfE3aq
+kCVBWzf+N8S8ms6oscn0QacfmpefvhTFn+I8A29Bwri95iNIQWKKBsKyYb/hRLDIhvKwyWH9UWT
j41ffJXiELX47AmUk4ouAR+9weeWc4wCnhckL3LW8GUBe3pPGQz0tAk1JNAz5Bv/E9+7oqZnR+C6
mL7jDOCrSfF3t7uov7GjEy371ndlwvzBN3QwsCmX8zpgtLhwAbDtgMMkA01auNrhsFG+okevG0Xi
Bk87ES++7teU0lUcmbZBSnZpIWlKfQ8kPCYiiyPTjWFM3rJjoR3ZHy/YtSELHEx1BCc9DGcGCKBS
35vOCU/xAWBR9xRSW+087mEc/fQJms0c2k+7Z9ZXKbeFAtYpDDLg7UH16Cb9N9EwQ1qzu0uzGM21
KUCI8WxwYeNKB5jBrsccN4Pyw5Z2PRYTHw/IANV7lSyt2t39UQL8xEn/H/i9jBce/f8gv538YXJY
/4iRUKAHdXzZ24xLyXgx69V/kcaSWlEdmQk3ce0dxpsCoB+CS7/uhZ7MfaBu2VyqzexMiQu1JyRJ
WeZOEPkpJuL4uAWjPBfd7Q0hud6dWjjc2wnBwXNWZ9Q7Egrm/Mzz2x13dCXw7cDdZO9IoEUUezjw
E5WnZ1GnjLtI8Vtm3Z6C4ICVwVkhPAKF07uBcrnHkgvM3SkmNZ2XaU4EWbCEickJcIjXb3Nnay2p
pLhKz5aBpBslswZTRkzkY+a58424xAmLwJIj7fYUg1v2oDZGeYhd8FO0xybD2U9qFTxMWon7N6gK
Jz60LYZXCFaCWjiVRABA6l8E0inMPmjFyYrmyVf11+ieUV/1suWO9YxhdwWEtmfnxmBJx4OMgjo4
uQocDfExFGw5H3V1S3JLIp1fmRcLSxZPfttxX/dBLDuVHmnWYk5xEwVANbbmypfvKYXpWOsnLTFi
LhJWAoQhyK0/Z670D7ATJ6EpPw4FsiRXDPkKytc5qIW5OD3IBGYVQAZ3w4/IEl/LuIqZ28tEpOf6
akMHNC9mBPmr2TbJY0S3Y99oHLomxN+NAUnQn1IG/fpH4dq/jgkUtUM9JifM8TCU99uT5VxJNnOv
gfZpX2y3xWym5cK3PDsGIRbYUyLwFYa9CVvoOMoTtMJGi9ZcIGgSF//DjF5GVPJJsNV+v/X/hf5F
LkRdiNGQ+OiPS+P0C4zqu5gm36ppLqS1ut3tw08167vgr2nMLk6fVOZxVXDHNpJDFOtuVkFOaS9r
gMY7KDvP705ubmMIULe5rl1Kiuso2E1pn4gFzhpQ3ft3HJ5yERCa3hfewITxq0ZHUa/KxBJ7uPKK
1ONzLH7iDdGiSoVfPpqHn+GTXTnp0lB0f8zEHG2Gl+shqrgOmjkswt0nlwdyjFTiNaVewjyd7aLv
ARl2zSlslFggjBkWGVacLv3yWRjN2fWutgHOT18fUBiMHSC5aZvo9mehx9ec8EO0jBEy2h/E2WNo
q09GMWB1kTcvjCbNYi8i+FC0CspBr/9uZB4QTfEWFnqdmGArtIDwWnqhlL+kxjvgQ4LdSuAAzfia
zdKi3SMEbzfFZ42JnU01Qciw4iU898LiAGFunaO4vR0E+AldpUvgLx4qhrbQoDZPYVdJojWmlI4K
hRWXBNY/wODT9l7GAt8cH2a7vXEbQHpZcCSAuNFYKLJY5tHOttEWFuMwwuGfevPyscrsclYVxQn4
Ax3/sRBk3THZd7xNIgA4NcHSjOOkMz7q5O00FQE6ec819NusbL/hXku645W0dhWEpQmtgPK9S0sQ
jp1C/vDGdZmc9RJB/bMNa94yMQSxH8XVn1yWsTwO5g9jv+jktV4V4VMmHzdrjXtDkfeOgL/mAjqB
DADq5p02eiILhLMyA3QrF8Mfa2KBeE0uh1aRIi6UgxcO3xRIV4BgLc0KVi51oGw6H8HBseg6blSb
8+HBiIK+B+ewcP6bcdE4wTRvD+nVqHIK85PgCtIs08WF57f/K4+XDidLjQ/e4x3RfTF8q3tUQkj1
822Jz4ZDs6Jfv3zSR92VWEn6fGx8Ju+8orm8xQMbJrHTDzpgm3UI+Rz9Mn2Jy/QRturyL7m30uzm
HUdbcASkV/ddbKNndZQHaPHF+/YUjojqTuvbMsZPXcCoaA4h8P0SUL0ydoK1jgs7daNBi9v5MTyu
URE5fJrITOIyjmKdSTLVX6WOtvyIqBURHiSYBqZrB7x4Isq/6uhc+7wOYm6MrmjocaF1CgOuKlt8
nedq+O5AxaNjotiB/ej1BR+Q+CRB2vjEMfB1Y7d/WcfWAWtrA6vnLK/OZKOv5AAQXdLj9cmKxIjK
kPBOCLmAdYZ9oDjgpTYFKIsPJ+dW1mZRTh9SIMfFCcO7K6KJY82UGtgcZ1BOoiAGmqMcWSx3ewtZ
xyjEeR9QnEzTDFWPrjwfpwUxYJpH3moI99QZdgRN2ZD/JVoZH+0ONMX8BO5swRK3ijCBnq695wK7
grBFjXwa4TgQWaNmY6F1tQeD0RtUtXGYtuZMa63K3u6gB/+bjr0PXQMSe0gUoh0+5kidD2rsDRok
4qWEM80zGFhLFw4MftnIPmsEOvMsM0BQw8fp9nGfVGjqpejx2LdhA3RPyK6cahfjZLBDIOBEy9Gm
5cLcDXBzUnGbfBMtYFPp4eA+D1Ugk0vP70kvA9OMpmVseW9E1jNUTIqAI2QfnHEVLQUQqtcjF4WK
zwuZ6Kqba42zz1y0jYiRSyE2SrG+2gfPbiIJsJ1wSboDmatNeFNMPFtjNsmUJqZZzqNfkZw0mj2r
STtLATGcDNWNYfx3HFcyMp/eqh3EGujIEiZ2MupCRN9qq54dAqXDfDvbl/jL0fNGPdxF6n91lpdP
AOI48pSNZhK3v/0t2g0LtG2GEC2ZuSBm/LYFrGoZK+U9MONg8Platwa6vlj3MGMbalyAen+1D57j
nBXv4WAkfjYtQ2/mrnD4U5U8RgGbydGe2ogvmr41w9wlqewLYbxh678PAJ0xUFMhUp/KaP3WYrbA
dhVTkWb9Sf61O8pWZNyyzVwAEM7RqOWG3F4ZZM+KFnKyTS1tYRqMel2GLDmpMxpoiBI7NNpCpfdC
fkEV9p+8V36sq3UjawjdG47ATnWBPYnBNPywAuZxI1IsFGH10slU9+2kUzvWiWP+dREV749puRtF
zUg72+IJC81WhYSnK8DhRi4m+pMvE+qKSgRWvK0PgME9MADHVGU2NF7vKtwaC1JArhLW0TU/Af4c
8tZDmClR5oOdw9L0J4AgeOBv3xZM8yaQXZvvxrleaUBJvTfq6Hd08My/4s+H7xAiv5PpsyLsNvJj
8P12fcff9lYecVg2XpamAynLP5FZ+o34e+mkGDM+5Ze3XVev3eLUW7VNqUBWfojyCHr62s1dt8G/
cb2uoDXnaB/ZHE+xBUWiwtl1Xdw+tkDFOYF6oFtXMtWbeIiJZ4VSsiWn3R30tRFJdmB9p/yWtwdR
vlk/CJ1uHhywI890qV3GZcKvkzisRPK9tSZO8pmSHh8JBNZptEPOO/6V8Iewr5xNPqBJX8+RmEpn
2SQo/gfnYNswEfwFML8Sa0FuZxHADzceaLWJsBCEsICi1iD8nSZn0e4m5dxX4kS1bgiAEFg7x1eN
z4MsEOQ+z23xpLu0Neiy+zEFCArY/k828KvQG99E9iyK0bAgS8oUU28F6zO5HVjjeiw7QJe6IBxZ
ICh5cIsZ7vmDBkTjpWR3f2x5/P5sU9dCtuw0DoHD3csiUW/lQa1NK3pSG7jSxIzroK9BA1ZyvMBu
PD3Aam+OfKelk4DCoVr/A791KcFrfwPWXbk57oNKItGHmyT0GwI0J67yGgpsSAndnsmXPiIIjPPc
eTyLyCXTOVZd9uBifPB9CD8q+dJBdEkFwG0qd4kBsuZoZpF5SR7ihBSqg+ZOCYEzRb6AYVTQlnbK
paTJyunGltoooyMi1sY1JP5C0HdxJZLJAxsrkfqzqZ0rVZr3VfzcmSJSf8l6lTTSEcuybiLS7P9Y
acBrYDe+8V/dm1I7tQYyMYx2tKR7HmDnIbQdUXjWdOcYHw3i4KDM7CA0QjpXdhmzRQgLd9PsVP6K
Z2ZksMBtiyp3puEyVSplPfO4BvGxYbA7Oi2USfSy1YR7sIycC1fWtsUS/YUPwgS+5Sfw6I/p1Cek
LOghzckseYCAMZpmh0pfT/tz8q4vNKp813/c5x0YvpBKtjBV1l9iKtCMHzX6cQJCT1ONKiQjuoYI
0N9GR/4tmdCypHwI/tCcWFTifIhn1c0UUDZir0RqlSakp2cKWkA3b9WKWc2JI834tjEd2FQYHygJ
ivvhN3JvTDip0k0GfmVI5/RVex0s+/LGQ5JYZMsajYLNOEHMhDpcWY2Ap5QKVNK1VzTFqoDHu8d/
OO+uA86++85jmlzz5MG16DpwcqIr9iDwSVi3NMZlev8jtQ/sRJsjMdTehz0Kq5KHsUnfzlcCSTZ4
OCwbxwn+9P1V3TLyBJZgRfSPzjvH+z72hRVSR21xWdUogyvOomjzjb6kTIGc4BkM5XxC+tultAtT
ZlzdNo3o5PoBJHbMGaPDjRzCpWMMKSLfmXdZwGTTgpt1WCAzvPlEfYRr6apSzMDXbchAvdpoNscl
WMYJGTaY0O7Bx4lG0gJdCo1XtUuaqHQHymwj+U/EjPr8OQSLs67fckN1soeW0e+z1UM9iRtqBt5h
KhriDK6OGWOUkwVHkrfut00qMzWbvAO/6PX/9ZMupnllN8j6z/UyMWKB1C9ewbHtoluVsAtSarvp
GSuzlF0PxLS8NnECgf7s3bXvLhF7jDviPjjt7PJRfkOR9bsdnoNLnC5mALlw0BBndxT393NV+cQz
P/g9LaCrliNCCXkgB+xpS2Vp+62Zl019wqXlY9J19Tx00Gbapr96okqT73B+2OcOZmtc7OFl6ekF
ijAJ9DC82BTUgA1pJXWw5U7qri7UOILsjDa6fsMm08oMtvBaa8QM5ZM2T2iA+6Lx+hxZmQK95cv3
XyR0gqGiA2S9SkBGqY9s8VjkpSKMnki8qYN7c+jR3UZpzM/QMk6amy4uJjXrChrQ9QIenAd0LN4J
C7mDOhZdv0kv4gOA/m3M7JW9UryvD3aV+g==
`protect end_protected
