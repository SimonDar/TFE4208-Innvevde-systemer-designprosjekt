��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�}{���cO�ݧ�Z�����_�Oȷ���-F`i���?nk2�58�+���%�9�t�ږS%���F(�`g�@>m�&�[ߪfB8G|wx���4�f�C�d�F��t��oۂ���G�y���N];�@�n�Z�Y�&E��RSpԞ�����	f��#M�+�b�����o�T���KD�J�i<ξ�M�������Z#�D{UbG���d;��L;Ƶ.�c����i$��x�(c��л7�ID�U�܃���� ���I�
H��U�1L�@����JS�!AḰ5�0��PܰAҒT��1��[1&T��U&���hGiSjK�q����Y�Uatl<�_宖`U�د ҕ�3/��nw�2���L�f�h�.�}���L�s�����.irhs��P��Ǚ�Kj�җ+m�t߽���"�Ζ�PB��H`a��I��lX,/w���D�td����'�[��(�H5�����Ab�h���\��	R#0R�����m@�WCG���v�� �x�ׇ��(�`��w��N�?TԘi���ms�.}�Yf����"5�����	p"��#�m���˩<����(gYܩT��d�
���K�?�C�*27���0����Λ�uY�#>�α@M���	�M-˸˻��=�(�Mf�AW�g��1�����#�O��/٤��Κ�;9��Ю�N��ߐ��E�l4���O�Z=�,d�:���Mya�[�oӏ|�B�������s��g$�fV������0������4���=:���B+	��j ͘�. �K����N���(7���2N�-��I���	�dW��1�K��q=��][���'H]�Ě�]��_��2 G�ד��\���v߭��¸�H1N�3�'j�X�G�3�w��d�]R%�!nm�J�Ʃ��^���5��^H��9߹�����Y���,_�{�4��:Q���FĦ���:i�9Wb^�L�n�%�lvs�oԺc7�2�=��jz��V�a���e*h�K�u�;�s�+���7������ύqg@��z����*�Z�*r���Ҏ���I���Ǎ��������a��G�U]��� ;��v(K�E�Z$޹؜��F6m���>ةI�&�����������X"ɵL��4)��=��t%�����@��=p�i��ɴ��2k��-�L��80��ǴߌX\�H�0���w�a3Έ�N��A/�3�$��hC��+�?��J)3�.��u!)D �A;Z�Q�[.���t
c��:bM�<
]TU�%]R5iV���Ґ��ǰ���($��SI���шV��jD��_*#Uo�{�F��ć�|�܆��ܜ���!���"G5	|._�
��Q�u�\�a^�C���]��"�̑2Q`��ΥB���o��>P��1pM��LB���Ǝ�H��.V�B��t��O+*���)�x�f\�H��8�L�,DJ���Gb0�~#<�[�߽����D{��7�z�57l쟩����Ne�{0���'���e}�)/�o#u���p"�b�:"	�o�1����(�{(�Y�)�	�;��^]�$���x��Q<������z����'P�I|Tu�aә��8e�yA�H��C�B�%hȰm��p�D��j�i����M�!!���?�n�u��p԰m����9Y���Ĥ�bT��-�i2=r%q��3�֟��%�9������yv6\��	\H�����;��������:c6I@��d]0��]a��W�#|� �o�����4P�?�ϱ��;�6�TW��$�F^�8��3�k�� ��Y7.nv���1c}F����%+��SЊ�	�F�B��h�-voꅢ�=D�+�#�pG�<��w�!�0�
�e�+V"�pn�|���pt#�]"�e\��uq��L\ޭ���[�)A���#ã߀}HWEy�4�8ǈhH�,���v����x�3R�q��Q:���L���A<������8"F� � �~�qmel�t�V��$;��γ�Zm*Ʊ:}�����0�Oq3{�)HI�D�3?P{9:�}O�e�>�\ц%|:�L�8��#3���F�׽�~�U%�4�<i�[���	,ts���lȬj�K���4V�`�	������J�=��؎g�XXr!��X�D1�j��=&|���}2��L�]vy����N��]n ^����)QP;I�:Y�d[���+cI�o�ن���/)�
@�=P����`6��>�SX��3�������[4�.]�M�t�D��2}�_��Kj�p��b�g~ 萖ɴ�Gw�s�L��L�v�4-�ǜէ�V�Q"�KήG�:��(�'��e�C"�^�63��c ��I����ġzb>�룞jT��$�s[�*��P��T�J��wۣ�' _
��n�(F]s5ot�d���TP�bvӸ���{��S�I�	M���	?����2=��f>��&����͆O�@((ޘ�0fE-s�N,,%Pyƴ����j�����4N�t
��qn,:
�1��ߪr�L�=^�	�O���/�D�J���h�tŬ�p�	��1G�����3�LN~��h���� ��N�W����i�u^�R�:X�	HV{흒+i���L��I7tp+��ϒ�-+��:� �i�vE�U�.}UP�i_�VRJ����(�����Օk��LZ�V��c�U�� ���3S^_���v���� A��̒V��D�$GZq Z�W�o5z�I��UV̇�>Ş��C����2^ �=6ၼb���)!6�G�o�M�A'P.S:���^������&B�u��|��m䑷�m�"6;_@N�Kde��P��_��>�
8� �Us��_e�Gڒ�\�@���T��Ju0��!"�o�Ax�6�0�4L��L�'�O��y$��Y�7��L��t�~B�9�v�W��yX���0F�)H�$��x�IJ��b�3&��_��i�{I�G�k^ߖz�.��l.�[�p���4u�	`h���߭��3^+�eq�b#�@a0�@�.bOשY�`K*�����1�D� 6���^A��"ڲ/���%���P!c�WZ��#ZQ�}��H�7�	�e�����X��q�����ZP��xnS ʋc�i.u�Qimp�s����A��,�K�.�(	ɚ(v����J/���VT��m�.s�:���i|)�����]nE�S������3���Ħ!�_��άQg�X����<�3.픦lH^�˿�r�ʕϘW�,�n(���u�Ȉ4|zay=�9N��D���MX�������lԨ�D福�ۍ�$�������B��*]�P�iB@?oF��]�	����Y���M��\�M= �K�[�H��~E1$N����&���H�8�C��El��kũSN��1BB3+f�k�@�*`��<I�`U!��n��c�I���.��EM�姘a���'�/�^O���t�Yᦁ�!�����aaz�U����fY���&G���q��n�6R1�C���(�v�h��7%�K~��Xy��&1���΁D���C���@��!�d,�Ȫ�`9�Ź8�)�D!!&���-�-PEm�\�`0�QjV�!�2�����uP;cl{��a	�0�U��|��p�-�/
�3ضAO�LMX�w��g8"�hu�p7_9��@z-�m&��+sM	��\�N�5�@vM��)���6թ��g8�m�*f�!��Et�t,���Jp�VνN��
�/!���c���l�c4�:(y9[���ΐ��0��LQu�6</�/�9�z�����bTGX퇲��Ug�w�H����yXqP�	E��J�Eitf��m`{�R����#������7�&�2�
?�y�A+@�64�*>t�[���R&���}3l���N�N�J������Tߓ�S�ՑIF�[׭�����K��v�����m\�\>�����P쟣z���G���|�^-�!4��K��3a.�����:����M�[D�+�t��4����'�d=>�`�0���`�jU�`����6�@\��#�Fe �`���f��.�T������74���C˓9�uE9���BM��u��6%ig���S��[�R�@`uԈ�݉~�f��	��|v���:����ɻg0L���6q�=ݒ�ʔ��#˓R��1�j=���3������2��>�{gz_}s)l�3,�T��L�"�EN�kٜ
E�A�R�H�(���q4�C3K}�S���@.H��PR^j�&Qx1�=P9=W��_����%�]
����y�<h3v��@���}�A��>��<$�t ��n�8�}��+�����a��c �$�/�y7����&!W{>�,�0%�T����̿��E�̇J.<�e�S���;s�F`G�OV[�)�P���Y7�$�T��F�L�ݠ�o�P��'��Nt��Ƭ��U����F��8�迦�U���,��:ĸc]��6���ڮέ��_O�|v���.��۳�,B�T����lL���W���m\�>�K�W4�_l�B�$�TT�N.�?�	��<R����q�����;g}�C�l�k7�;j�Z��<*8�e�LȦ��W
Ο�;�:e� �Ν9Yo0����xzb���ƃޒ�J�]�M�(�Z k��S� �#'υ.��$Xd��s��:�yA҆�J��y��L���֍�d1_"[�j��]��Yi�	��p�[[o[e���3e��|��ц!�m����Y��&�7�¸.{{�X� 	�� :�w�5�,���c=�т���iI���~����E��sڷ�~'{
�(�j䃘�ˍ���!������Yu�~��Y	g���M�(�Q�L^��9.sy�lR��yݎ?נ��u�e3xS���x��!�y�S���ч�R�����Pw�*n�k�rYKFEGQ�1�-�;�ݝ�<O��nHo�C]�8��q1B
��}���-��4-�d<�� ��C��`]�2�Ѵ9/�����i���G5�{.��[��F,�JE�%a��S��0Q�e�zT < X��/M��6S�zYޕ���v�[��d>�ɴFP�C������,��R�67+�8�AY#������&���Z[ԓ�O�P~u.ЩC�<���.[�A����q����bh��N�>�m\�1�;H>9*���Վ��-�.q�s�������['��OqȦ��oA�j��҂�|v�U��<��I�����.��Ac	����I�2}��w)�w/S̀1ri�`�	]�I?i	i��I��mw��y_� �l�Fn����OO� }%�Mab�Fú�E�П^፵a'�.${����Yهo~7��1eY_����6��! ��d�yM�/}p�����bN��8�@���҅�x��-X1��7���P���xw~�F=�����idq��?tZ��BFNG#��"6�$]�]��7���Qr�i b�Ԍ�%����G�[��������3���tq��cPU.y�c����S�l�y#,_�8�3��b�_ +��ƨ`��B˥���S�|	�  ��L�q���R�,ﻌ��Z��W���91k�!EJ͟�[P-FW�������@�/sp��h��YeE��Ыi��e7�S�c�&Uѱ4LE���$yđ�㢯�E]����B�|-�ර����kќo�G��Rc�[�@����6��&���#�j0`�=�7f�Z�����"�AӈU�r�i+�ة��Ty؅ZIm�g+z;���S�:"i^;��L�=ς����,hB:���l��:���F����B�c���%���Uwl�[Xa.zYi.��'���!�_B54(�� �?*�u]�����\i�j��uz��W_��5�x!�������R"�܎Z�ͽlc}�JM��<���4h�^d���
���i�J����E48�3 ��6�T����X��v��,M{0���|���Cb ��}=?���;�����ޟF�F�B�C�r̎AH,%c�3|u�ND0S�ʂ9�����vмN�=Vo�C'��|+��U��[���֛1P��}��i{Z����a�>�<8��@.�iṽ���?�^���DR_��aH�>A��P�/�����yaPI9I����ކ�m�G��qa|Y"��C"2�~�St��댽��_/�UfU�pr�"����uy0ov61`֕�������ݍ&�@����-g%���6��H¢������%�1���dL�j�>)r3T�k'�6�r����dok3��^��ª�fӕq	9��bs����#������6T_�j[����I����\{և�]��0|�W�e� L6�Y�|�J����J�-ֲ>A]��!�k�IV�/���
��t�Ñ��6�~����hq����?^W�Q�V�(~*r$�z�Pd�r���Q��
އ"�kO�\'!�L5��=,V`��ґ_Q����.�6����m"�s�+�����䝗���U-���w`r�S�UqeI��I�5�0��q���˰�Ͻ��2�N�fJr�C��� ���c�����WK���K��~	�Qx��6����r�JD/;��?�7��4��@dp|�V�%�b�J�1�qbwUA�
S��,��!�b�7,�2�4c�D+��1<�p^�{�T��[?"�.z�dm��AUf�}��W�7ٙ�/�ѐ����1p���K~V�Õ
֎��jq���B���eǮ���x^]RQ_�uO��iZ��}[K]w޽K��J1�)t$,Y�D��ڔ⮌ 
����J�2�V����-[��nY�nu�fɇ��t����bS���������Ī�h�%�g)q�ݶ���9:���U��/C'� k�[zf���$�T���8��U%�`���c{�U�\�0f�v8WM�6�;]��ࢲ��߿�����)/o���n��]�T�8�s֊��a����[z>@Jk��2�6?קl;�7UN���Ѵm�:
p���=�y�I��7ۖ���,��4�;)l�p���[<�Vr#[.�^9�d�B��'��®!�� ��8�^uo�:T��4�su�ņ'���u�
E�S����GR�� �<7+Ѯ޸<	y����̾�>c�f��˛R��H�g�I����,h+[�
]l����Ϥ��,��������My�	�]�x\�v.�@�&��,�o�[�(�r[�����UT�s�4E��T�"W���B�G�0��/y���{�0
%nq���ЬB%���wy��-�"�V���&>����X�^�+��
�#�S�㑟��L�����*��Q����q�be��=,�l5��)e?�1Q�ߥ4��U!}�!أ7�KcDn�q*��3�֍�g{��o��9e҂(�n�!^E{"����Hk�̣f��B�`�	`�u��q �-�V�������}����n=�jgY�u����N����
�=63_K�y�=Ԋ��<��Z�	��C+��K�n��a�="����'(�� �j�1����Z�PIw'S���咙���euC��\!��|�ZJ%�LTC/]#�+��������R�kZn��<[zC�$ڛI3� �,L��������MN�� �hN�t�0�����"lb-~WU%�gg�z|1��<�CzcN��~��cq�;j�+��o����(�� ���b�ف�,de�^nbz�}�Zr�]p�-�;�$�wϓi���9Y�_�B���`y9eL�lק�Uݕ�r�`�	��1�k��at\ȋz0#�th)1l���S�?R,7��j�&��z��{��=8^����d�X�mH7����`�e������R~��^�J4�� ��Ñ�-�s9ix�a�X�@n��90ܰ.fc�G&�=L��0���b��u��8� �l��J+�L&��ݯ��3�͗a2�7��R3� ����&=L�X���/���N�k���!���9B�o�e�l��w��fQ(M�C~0��2�&��7TMD(k�er6�[�O�A�y������_���T�	�,ǁ�׏`�����88�ͥBH��D�?$�	c\�t]����`2
"N��������"y���|�^)���)�5�H'�"w$s�ɒx/ߔo?�)�(�8/6��e``���M}����Ӎ���`0������H�̛�-��Ԁ7Q�������5�[��~�>���C��gln;�)�u��}�/�u��hC���C����6Xf2��Y�`�~,���#�1�TSM<.�m���<$23͒ ��d9���At�N႔2y���j|	Z�I��@��<�����6�������L�X�}��L�m̖Z�˧o�*/��W�B�<	�6��)��
��#2��@BU.��v;�N�����_�I�:�*�Ŕ=�^�_��#�򢩛�������G�e�����D�S��cX�8	�����L� �x%��5����`c�7@xq���%���漴�v�_�(O�V�3�H{�̃�BZș9��U���w��6c(f�	� }���c1����+�Z4!�ɿ�F0���?I���������Z0��T��>��W�})�Q��T����~~o{��m��LZ�a���V`\�)d6�������G���H|FS�d�l8J�Y�>a@NrB%��V�d��	��|��C���9��'m���l�T>6�nĬ0{f�C����LW�Eo�SACpK��q�='m��͇8^��V/�[\ @�H~M��X�=�Kܔ?��+@�/¡�M|�ʵqA*9�������v���?��GII�����=Z�,��F�;Y��a��Jl��-��s�
�Z &��~�+�[��Ɏ���K��;����'6}Ə{��� �������T�E1�͢�����\]�)�_��8Y��Gr%���7���"GbsoL�z�,����s�W�Y�mR�N��r����Ҁ��R�t���r������08�['"����G uh�������Ǆ���	׷<�{h�"��Pũ�f^��Q��$�����t����t���/F�w�.�>�+P�� }��?���厓�f�c.�ng��\�~!�i��SU�q�鮯9�}W
�����3гcd?�ovQ��F��id��7���]����K���XA^Ov9K�ܝր �xd�?ܼ^�@a}�%�s�-!Q)@S�rh�HO�\w���[Vmc��&E�W��0��|�x�)Y���+m�J7�$L�z�I �J�S1�3���z
�F�&>��0;RhUh:��P?}�KD΂%ɖ0·�Q\*�BP-ZM�����vgF˅��D����$��xݾ�f�l�S�iaK��������c��g=�v5��$������O��%*MSג�je��sܣh>��㨔��E�t����J8e�0lc�L�:~���Ɔ�833C����3p+ŴɕH�]�ų���cBׂ���y/P�%��N'�72���'3?mnC��
�D�_Z�K��J��g��\g{$ݬ/�7O?�-Md�Y9p�p̭��X�<�`NXG,G��=b�rȌE�9�B�[��~��6�&7��s+{*R��Z_�[cs<��4D�S{��Q-��<_�Y��"���c�J�Y0'w<���Gp\M�~�,�����F�\�-�/2��K�\a�h�$0«+K@L�]�½�ԓ	XtcNs�S����>(		F��Whŝ|T��\S1ZR����i����&�سA������'jX4P�Lt�B~��Tj1M+�L@Y�j1E�B</����r��i]���֟����R�q-����!�	/9�;�4�!`��
��R(2�1��cW0+����꿻���:�m5��X�1r9�>�g�<!��d��T�Qڤ�p�n����Axg�
�R�1GV�N�}�E�[s]��$�­���'>��k�ҍ��8��6,���0�+���b_$�-�L�Њb��͹�3ګg�-��?��|�_�N��l���z� $z�}�� �r�X,R1�F������R`���
VR��\̦=HTvY��⦧�W5F"��oפ=�Ō�<]pdz3t:�D���o���_�T�~�6	�H�7�0�n釹���&���/����7��?_G�n�����J���R<�I#�����U[ƨ�jaLlb:�OCۮ~'WZM�:��p�|Sj��UR�[�U�vTcW����!@��<u"9�n/\k��I��W��M �ZS�WG����<)�u�Z�]���H�-�Z�DL��k\Tf��A��f�R�n$�+o榆o_0���?6m�䄙��H��.Gc�j�F ��t�Ҩ�ۋ8"=��G�B�n�7��ڱm�#��7���q�z�P^�%2c�e�"#J�f
)�A�m��%������-�/=fy�,��z=Z���x�r���O�L�Hz�V2���	0T��������w8�ji��VX�:���ih�F�:��ś��~J�&Ŝ�v.�$�L;cEV���ݘi��X�h�Hi�z�`�0�҈[e�"��S�|4_[��ja�Hp~���v�8�I.��R�܇Z��V��֞�E����숙����m����Hw�i���OKl�`ͬN�&�k��k�� ����Q�|���N����t�A
(qw�@�쑶�(�V��$�ă-��$ �%�j���Q�X��)�*���jW��(��0��Mp�?�E��~E��xDX%�$������r�e.�E�&����>��$p�Mdہ�VW4�dM�:O�;�\H�[�&L&}RؗQ���AF�<�xAy��3	������LZ�N���ڬ��p�z��q�j��a�5.ȁ�Oo�@�4j�����-�d�tG��������(������������� ��ݭ��^��������?�^�I��'��lY	]PZZ�^�z�۸f��	��e���a)[[/).$Ҟ���'��L��y+͝���%?5�ad���Њfd幀?t�m)?Tv�oz��rHȋ��Ng�n\�j��9�#}����pH�$g�bp� �7��%�"�;���j1��Qh��"�c�{��4���.6b󯷺_ŢG싍����x0(%M%�"��">;�M��N	t��~�f@{!fϸ:�"]�X#�M+���5�Y=�d�2��v��E�,ێm��k}x�γ�LG���ʁ s+,=g_p��bZ�DF���<ظ��zZhZ��<�5��]�G�ce�W�YT���:�/�&��3�����l��<��o���E�|Dx\nZp�C���1t,���� E{b%V �	�3Ltcݤ���?�V-�^z^߼Z�hD:	V���VV�?h1Ue�7Q��G�(Z!䇺�Eߚ�\����L�|O�k�������+��d�'�y%��Eq(Ƿ4bJ��}M��i��ȵ�􈰝&|��1�]�O�&�މճs�d8\�s���'G�1�(m{��m�H@"�e���s������>�hi@0d �A��^��I`m�pP��5x ��lV����T�Z��mr�+���/�6�$�ڰ�${x H<l�7�R�z�F�E5R��/�L.�U��ɬ�5���2��D�۵z��s���x\���z2d���~��=a{#n��{�5EIϻb~�Z5�	*��T����� p'�2丢o,��O���t�������) Ǥ��&�zD��� @K"ԡ����̄��Ȗl�p�mf F|.�Nal�8l�>pr�>���;Br$[��Ήy3���{���ʼ�A,�1P��Fܮ��*U�VR
��r�BE�|8�O��2 ���=�v@"&^[AVH���[n�chv�D��+�?2�-W�%�7Ř�ܜ�֢0����\Q��
7)}��t;��P�(7u�����ci��@��m(���sFQפ�Y���2ZΞǕj�Kw&�e���ֹ��O���:���rFsː�y�<�jzSC��xm� h��F���/%��y��U��i'� 씕���؟��Ҷ�������u�[ �����{�~�A"��=�=���D��HG%'�rEP�N/�X_�e�A�ul��(g�b�����/9z�+�t�1��L�?�86R��7�cX�w�����,�t��+'-���?���|�tp��'0%2e��/���[�2�}՘^��M\�̌Z0�1�t)�x:<e��g�7N�Cis3}��?ٛ%�O���~�<,qm��˗|:c��X9:��Z� ���8��ļĘ�%�CB��u!6�����^U��A�� ,o������^/Z1����O���L[b���D���:. ���� ���n|9w��T�=��OO�?(na�13�ǃ_��̚������adq�������m`��(��M�;��E�*�����o�$,��OW�X��W�zA�c�O���N�6��T�����730��H�ԧ�udn�Ѧ���ϙ��͒_8�@T�w������*>e�:�{JE�نꈜG%͞���	n'.���t�.�C�y�<(�\�`ޒA�]+s�����^0���\�<)5���N�R�y(���3C�I��Q	�kQ{���V�l��nx��oI!�)�Q���J2i��L�e�!x+�_�"��pC[^ _����G���w�h�e�/7�OL�7ȎX�f=U{��G���a&�����PPv@��}�y���]�U@�y;d�S$������K�9i��`���w���1��G`}�GIL��O��O���s/�2#p���7+��U�+��j�����E<��T �5E]�d���`m�#{8j2�V�����G�q�dLK>�

�������eF*��z���c��P��:iW�Э~W��w�?��I�i#d�HL�|�~�� jw����H8�)�bM�w��p�� �T���SD���@��J�@
����P�n�Z�S,��]$G>Y��Z�7��/���f�l�@���$��sy�P!Qq｣-"ky��6;��W�I�9�1��sNg�~��gq���E0�;Eu�����je��=pK 4p�.]��[5PzZ ͡_��c¬��f�bR�G���ƈ����o��F��J�MD2t���/õ�(18`��#�[S��C�a����Q1���
�ʕ�+l��(�,̲��Ԇ.��%(-rV�m����i[Fc��2J��O�c/�
�T=���m�Wu*���0�P/7t�z�U���Y$���^�t��v����P����F���EBE ���%]ZY��}aiK��v޻o��>'��AP����\���^XwhjsM��O|�����MT�) �F�	5�t«+��&4;�R����2�6y��m�/C%P�S 0ۙ�y��gh�.�'�I�;Q����y��Ķ�3葌OH���#���(YOlyԵ(�#��M,��[9��><Q��L�v�P�?w@|��U9��(�ay�Y���H�
����y�٨!��#���;��+�D���I�Y܈�n�|/:�)�Fv�W��){z�U]��w ��4D(-C��gb��3`�
�?���u���&�x�rމE7����E�C��%"�"g7�K�c�+U9�Ȧ�h*�(���'�S�FT��`���fI�Xi<�!4�~��Q:{ 哴�&/k��/�񢡳�}�"��t+C��[���_�9^#ĬSDh�]�L�
�rg������C	��
<����h0�ұ�s�*��Y�{ykPWD�4�a�?FK���t��$���>g��ț��|�NGc�Δ��:��q1򆶹��xn�,I;������?�X���Q���c  ��e�u�s0��U����@�!� �SH�\�a��E��$�E��J�;r�p�����͆�	�1������8i�MDp���������e�2���K	�
Ǡ�#��]�"F���Gf	����A@.V�����F���	��2�?��FCV5� ��&ۇ�=[�H%�d>M��6n��nh��L�W�':�q`�h���܉	���RA��V�'�V���	��b��i4��X�b�$e�	Z����.Ubbm�^�G���� '~e�ȟ��5��=v����Z�+u �mN��(	2굀�}�>�9��s�)A�ȳ��f��`�C�0�� !�_�sW9�3�L+:�UgT=oxuH
�qz�4�B����n.�Q)Y�n` �mC��78����7oZt#n���㬙s����W�� �?���8H��k(��_��a�����I�F���%(JV$+��Z8���C�X	������G19o�Si���Ye���O�;��S ��L�E����G\��5��.b�ML�k��i��)�"'tR��G�S'/zï�.��z��=H�����Į�D�q._s�N����.��OG�J������`
]M3���2��>�v�}�ԕ�ۘf�L$H����Q����XRX� ŅE.o9��2��D�{�t�7V�~����b�^��i���:�t�k��Wa�ݩ�'6�[����m�5�>g)����u�p��XZ��)B>5�S�]0\�k	���:�*	�p����ve�SX�^ʄC�����ųM	��d�]�e�"���=�Z{�������G#�-�K�.�∭Rni�+*��Ia�O�H1:Y�!���IhI�h�K�>��(������Ϝ�4ݗ�S	f�ϱ�j�?�(d�"o��}1X��)�5�F��<��m�`�YU1@�"�OS��=A�;���cM�9B��?>�O�{G|�W�U�����S�ܕ��҆C�N�P�)�갭 �Ǡ��U���:k@�|%u'��ϫr8�r�;&h�F�ǻW&L��&zn씈6�,IT���$C�r�zj[�=!}��b�&0�'�˦@V ��J�F44�d5��TXc1���>����r�)�)搦�.�X�l<M�P�2'��֑�Q�67������1-��"�Q���r�y��_|�����U��jH��5��g���I�����yW!%�x��6��������un#lXO]�&�nd������s���g.*@�^�Ձwyҍ��t�>YE�5'���U��80C���=jǒEޔ|��4�xbO������{���Q�B�~�o�)��@�`��cck�}���M��U�|z����y���/	E�z#�jP�.2�W/:t�PJ�0 �����s�i�d|;p��-AJ]�����I�������7��#��}OU�]��AQ�B56�峩sMժ���t]�� C��:8e%�<U+2�ġ�d�ܸR�mfc�|�4��e3"s����2�`�¨֟:��S������A�����>��Me��� �k�{�]=��|��7^8�jpg�����~.�?������i�Jp�$l���pل[f&���B]�v0��*U���[7]�fQ�N�^���A���r:ZC�'9R-2E�i�>�,���BT��d{%�N�� ���L��鲝C~$r0(6�$Q�6���VόK��]��)b�eT�
.����3��F
��k��fj9��jLU
���ْ��抿��76l���KgW�c�~�-]�έ�Rɳ�h5W�C{Iб�p�h�b���K 54�8��h�*)u��ai��b�l�v�[ޣF�`I�|�5<A�.~`�����؆p��(0���l��n'4A�@����֒����f�H�J�Б����k�\V;��ν�o�^�UDtR�W8��Mr�'���TUͭޏ
�j����E��%���9e�^.{�t/��MH�o�4ѥ�ɄL��Z�W��k�~�nd��r#��1x=.��YIs��������RQ\B��zs�뾽��z��i��M�[M�vڴLz�˛�^7�3�O��nen�_�v�*�k�1��S�4��v��Xx���LApơ��!���曆m������Awe��H_�aq�>��h2V����o�G`
��zI:��-��Y���k����.�4�0�5J$[�i5�w]L����A�k��U�fc�����wޝ�(j)�ՠ3v�<���_W�����Kjks�9֠l[����dX qp��!cM8�x����v]#����`gEx'�� u��vi|��$p��E�"�9O_�ʐZ�7�0;4K���n�Ұo���E.=Ѕ���xJ��z3�d�3:��{���[>xc��4r��n�:����I��/���D���T��3W(��l�u�	K�	�Ҙ׳EL���+�3����{![}�����)���Pd6SY��o��΁0^���U�M�UE��_�X֤��A�G��I	��T�wf{R����4�\M�l��>�终}z��@Ӯ+�MϮu1a�"�*K�j��N~�9� Ý���}�FK�����β&��Fӵz���_F��P�s)]P�͖J�������ݡF@z�\�@���L��a\o�Pڣ.�iB=4A�)^�=\����_������1��$�U�������BY����qD',Y��]7[�����I
w$�v��s]�$�+k�!�X��!���n**���GU��g��ùnq��-�Me���d�~�Ҥ��"��	��ט��<}5��7�g6��#-U3�-�ש��d2��U�y�͡�pV((�Fe,"۴��M@����/�,��̔�
�ֲ3���tT�/�����%�l���v`�eX�OǉߒsS6V)��q���pNe�&�^�p��i�99��9����O�P���ſ{~�<E�M���N��>,`ӹ"�SZ?kQr�pP���3L������;�,`��.si;DI�Ƥ�m�K�w=�����+Z�38pHl �>�&���=z�>g�}�Ӡ��Ӽ�`o$W6]��!7�&#m��'��2>��@^f"�>��uX��'�/&���18$I�(��Z[�=��s���(k���[��!:3�v�N�P.�5�J��?�x�|V@���ƥ1�b���/����#��N��,��	��8�)�խ�L��8~���%��#�����u���Mw�keM�s�0�����^�,N��(f�Fqʵь��?��g�T��7ˬj.-pi3:��a'p����D�}Ov2�\ޯ@����������f``�U>�@2���)*�� P�:��hꥳ����T=��A��5fd�����\+�6>�ka5;��\�//}�/U��m���Umz؀����y{���U��l��0�n�ן�EnE�)�>2�2t�����L��6J)�'g��	O�P�(�}��`8�a�N��@gD����09�@��9���&�!&8�y/�!]��rgB�2}E�E `1�*��;���oF��z�>Sg�P�]h2���j�����^KFt�4 S.^�kb�}��N��[B����,�̢!"��3���S�c!v[{��	b����rc�\�hH�4�/ ��t2� f�$-��s��JɑGҶ
��l�u2��~BF-x������.tt�x<xN��~��8����-z��QV� �OF�=��s�:��D����ѵ�ߏR:)�#�8�o����@�@�͋�0à���]� �|���l���S��Ѫ�JZ� �'�.��˃	�@�Ɓ�՚��:h|���������Ƚ�Fs����J�g�@���g�c<�iAH���������մ�^�檆K����_��Pi�]�LBhn<�#��/3��x ���.�:�����aHx�,�Ch���<pQ戦5B����������)L~D��7P��_�Ipс|�J���D�EA�UY|��fp?�w@��Ӄ*Q�i3�C'�X['����ey��Z#E��`����ky
��SB�`[�3�L���*�k����k˴{q/�����u6j��;M�r<��ٌ������O%Es!)B�u�wk���	����/n�X��	H��o
�ʸ����>֦������܇��F����<o�eʧ=���^�P�@��� w�F���bXl��0���� U����j̓	�^�%���p�@��E�J+��pW��m��o�'aQ�G�zb����[���PL��t�Yz��<� }h�2�ز�@�qrr_I��Z��>n����D]o�J9Lxb6��P[�g�G*_52Vv��Ww��I�Xw��a�����!w/l���3�!��Q��ZU�z� @K��+/ސ�[틀'�ݨp��c���F?��J���p���RӛR�jo�[��\<�y�}*\��z|�s�ۭ�$��p�������n��C�� ��N8E�-�	w����ۇȨ��V(�|��DgX�����������\Ho ���Zw6��q3	��u5��H��~��%Y���̧b�խ�9N�;���/�y��׬>	gC#�9�̲8�\��\z�K�����{�!�jg��J�xs��Ԧ����#�\������< �#����M��6� � �S��d�ǧ��w�<=�Y�⇐�@/�',)�٪Y��?���
�`��f���\ByX��v�B��rY�Ci�킊­P+��������� ѥ�hq���?�rE%��)c��.F�%��}C���y7 �y��BI���������#(�'G��[�\K��p�/`1#M�
L#�eu��T&�v���[=��������Ǐ�̻��H���_�FXY�*>�T}�q���
�3�/���	۩p�����vF�����#�
9+��7h󑡐��g<�N��=��Z.u�����p�N>���`'aCW\�Z�>��o�4V��Cm�������B�f&ʜ�Xg�۠�<�T:;���U�T��1?��s��#�g� �0r8\�,4O����R(o-cb���Y�� ���`M�.n9/��Id��?�D��P�f�H@usS�D��Xѐ�]_�!�7���<K-�b��[��M9.4����;	�ǣ�P���z(
�תп����'t�x�����(<nQ�S��7��i�K̾��.�L���|(�/v'�ب��Ҽ�����Y��GvP�%��Zۀ����Ѝ�X���<��+���l��o�T^���S�Ms�9�Y�`=���-{�%P헊 ��#Аi�>hz���K��]�vP���S� f��w+��������{�^:m�5�6'�j��d�˧@p��9V�(��������g]v�	Q��op�t�]��$TΉ>�w�;�9�c�}6!a� ��?�yOe߁T�������p��V����a+$�T�<�ZLi[��HqN������ʭ��T��М�ZT zyZi�,�M�dq¼�q�� �d��O0�j7��^���r�k�4X�O���}�B�0D"��H/~8v_��ƚ�(տ`�����������#��9���U�ìG�b���W\�C4҄�����jھ��}�[����+ǽǁ��lUZ���ar@D�LVÝ9�F{�ﬞ��|����f���~�O�0 �a+�Mk�>W]��iOɂE���� �*@�������WF.V��3�љ��a��~+/��f	L�g01:U��/1���P�h�q�A���X�. ��ȏP�waW��o�d4�47g��p�*̝�~D�2���!ce:�pչ?�Rį�^�ܲ}P!�M��!Wk�+�M��&��@8�q�*�"6���oD��0E]/�=ҵ���=���w�8����F;E����O���E��ѵӑ�F^�^����{�5���:�XuV_����w`-a����χ�8:�t؍����A���t���C?�ł\�uVʪ��]����2�.��wT7���R=����d�ؿ�w>4���/ӪvR��?���w��><@Gߒ V)sPSP`|쯃;Zo��gMP1��Ҿ��.����~��%��jl����9/�_J�x�z�f�G`=�ƞ�cv9��H�1����0{��_��w���E_�sŚ�u.�[�jʃ��Z=
����N6���V�O8���>2����n�F+8E&�g�aϊ��d;v�G%�?����O
!��!]��J%�'��%��<b%�{5���\�hB^�R��H�ڈեY���M�72g�0(\kV��>!<�(�a=�y3��,02'�β�`p�6nH�� c����v�}b=��cc�<+��'S
c.D!4�!Pl�m@q�R+�e̙k��:#�Kq�鹑��%�b�j]T��l���*y�xƳ�{/]���g�;��<[�5n�_�����֬�崫xk Ŗ�b�|F^0y����wT�J+v�~�(�5��2Je��Oȇ�&����q^f�B���f�:�rY[�49.�}��9~���;�y�ߒTU��?T�{�nȃ�G��Έx�M�0��F�|�>\1��yJB��y�6Ѭ@�7�TX=.�<��A����m��;�0���fʪй۵��jE��E��
�{�3@�
��f�_me��bfaB��C�v_Mb��]�Z���⓰��p��$Fdd��J�y�-�|��2��7���R�ݜ�$t���@2����o<�w
�J�a���vE�@@hj8�w�� �O��*�D��,��p<�07x��Rv#�_M]�<�dr�Q�� �3�����`���7s�]u�QRe�g�A�1d���e:��۶��F_�r��@{D��%�IZ5�~���?�5��5/wU�G'=��0Ѵ�/���U�hE -j=�:T��3���4��П]��^:���ӷ���R��&}�����}��0闤P���;��;Q���-��,�[|qbV���U<���R��/�/yQg���4(���:-��P F��o2>$	c����(���3N�04��F�u{x�!G�����I��2����D�-���p������y迠����9:��S��P���$CV`[�Ιi�,I�V���=i�qy����^m���+ ��àW^�k��\�E��V\�7[j��+�\�i�"�����U�ڀ��;A��m5�A�x>.�Re��;�]�'��Ɇ/C���jy���r4�˜����I����l�����	�$Ǵvh�;�Y'�)�K�NƆ2��
�+Wl���� ��Ϡ�E�{�2dp$1zb��;8��m���r!$�I�]���c����r`ӡ�򇍘R�Kc��Y�a��~���4WMm5�h�-�Y�I�tA)F~�F��~�){V8�ҧfm�8ӝC�T��Ո�M�Le��c