module fft_source_interface(clk);
	input clk;
endmodule	