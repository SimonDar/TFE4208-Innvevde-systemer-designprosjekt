-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pKaSCmYtZH2suc37uAw/LMPAeLVBXbMabZiCnjtJEmzMC8TverIIDhMiauA/44hA+AdEopxFWq/m
03bN53KxMuF3jNeEsnUg5yUphk2MEVkicQD/Q2ttVFwAvvAJmNuCmvA3jJkW3xkYKsp5R5eAR6Gv
vmilIFrcLp1htlorUy7vpZvXM1JQn2Tu2pN9E5u1ISzZlTYKrItgHF7mwt+i3ZS2EYL3I1SXvipB
fRh289HUXPUZkPgJcPIxdLcYyNmC8C9xy29hy9hk9AK7Y/GHVRIlEpnms1wd4BQHVPVuBel2w84i
OMH+tIF0XkMIkZE2gY9iqK/kCgqRrso7vN0GNw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
2Ip/ZiwxCauZXuoFO4r4atCZwMzRtsAaD7v01oDKuDSj5BQO2XTX2fRfHEx4XB9IGbOpep2+xfcV
n1bDYayBJK/AQjjnttCXBy1xYEhptarppZRkH+OEAxZ9gJXyu5pJ+csEdCob8pt1eiaIuvycgm7w
f5yo8IiudLQ5OPmLpvcXiUn+YKQtVR4WALACTW5tEI1PT8UjUQQ4oHT1MzBu3l5UAt2uze5+pQqG
0Ib+HWjXRTaNhJYwauMwkvnCbD2ajRK9TfZnw7/keJK250olnLVDQXy+MS+cYBb7SzQxdZcefEvT
k9to428es4z5weYwDN6avNmXFxfF1NmLwLe06bjF4NUn/zCinfp+UA9L0x5fRAjiVV8LjM64VIOi
wclNEZWslKxkgyUZvJxl7uokDRkl2cl0rYUfF4ghaaespQWbyOQPag5xAalvJOTRRk3NhrTTbJFy
uYCyv3L8Z0hsQuo0VGmYY+RO+JoqSFt3UN4e0ooAJJOjlkmjRKQYsEec79K+kZxlM4ov3mab9CNo
Nw3X2GlLbHFaiVvnEaPx6QfQhyP5mWjuTujxbUvz5b1LP9IFjthmfBS0Hll5lFoT2/FktRVP5K3y
zFtjeCQEW490DGSgki7V9L3+2yqovRmnFY+Z9mResShTjzfictmPJk47ZNJ/CvlUivdYTpCu0RE3
T/8B7LKEo381m2+zPNqIIxwc3BWTqZhiC9LFR2Cu6AFUwNw/a9p19BeVScmFtU5i90qCgtNUQuRD
vQYIrEpIG6l3edzybVakrFAeaK+0Sg2CqOa6CeBZ75T05K6OQba9S++/XD8b1NEoeZf51vBIV+2k
/+WLgGwJOIdp+TGW7Vdafzte4TbF2nZTSjGd9Psa32k1G5VygN4nh17yh9grWZ4o6sFPhRV5d4qi
ClUs4zG+Jg0QsYgROVkoZQQNp/6PKdeP2IxFIITJjUUSQfXkETCwiC9n1sdWZX9zB4fus9r2Clmh
hf3ZiZUIe51UW3gNjbZY5pjeWTj3NGSrhVK6NaWalOZmCENRQ4LTtuK0zkOw2A2x9ejJi4fnVGNt
4xYYjw2YvNVT2yKiFLe+O/NGaPxtuoEpw/zJKCS1S2TE3NJWpRwiYo36XK6tna/eYDCOWcPXzlC0
pjl+yloXTOZGM36g0z3bx6DBHxmpMlbdkgphtE8p3q0SpC8tncj5hBwGDm0sSzZbE2QXAMyLC9mo
0D3qDOO98M3Yd9po+GZ2vVW+3jpKisb8nBxTeEZ0rbA4uJ9F7wRp3B4AQLIAWQh6dohEscUKdBuL
MOJkY/IRz3FsjdYi6/TX+Wj0GkKq8ECFn8fkwANzU7mHtUvc0yJw+XfDYq72U6FvWu2EuzQgfqEG
cpZXrPesNe+Azo5ZC5M4Dz3R/sKyS0ZSTSz/rLPiBn3kKYi+7pKm9COt6l9e1cE90KfpOtg+iq/U
rrUQ5QkXSXb4YQ/VSTIV+FEKL5QKnk0JhJD0ydjNWXu3bYH1B4FfxfwGoNq2oEJ+a6MxmYLfS2d8
cgDm7eUcXekpPNaWfJ7pxdG2BvDVnI0ZOQKEWGtDid6kQa50cH8ev6a1oU+okcSpVbn4mCgaSLaU
mvbi2vYTUtiLDLQFDHd3xfa6WlVWbsOOiMp8bagTbHnC6SvyOzRyV1f4j9ynrmSHbLmVvWMGvdRo
d5Pb46NNHfLHVtmZjv3TLzx6FueJ+bPHSr/FQosMnLooGAYd7Ry/rI0Nqv2s9j2YEj+MH0BfxM2j
jx9gwXQroh+zVIFgmgu0hGr57s1lacz3ovGQ1m6iSJ3w2PL8bU8YwaaTvv0jltV9NR4TnrLNwJO0
h0M2eexLTKO/A15v9RFMlKXBOjIt7Xr0/FCRH38GJ8zRIBinmRwJvzh7NrazUmcMA96vgUmM/pV7
L0YNZ7m6S1izZije3VoujS6jBPk2RbnF4kpeSJwfDVbYCZhs6MwWhiP7jffgFjIYpuVWqg47MTiC
jowmnz75IEDkedM9UR6k1lIBUMZFqwagyZkEWKApLHqqyOHMXSxuFdclXT6aE/Wm3dJVnqIS2FvM
ws2tLjepIJ27cILV4i1Bim4wJDXCsK1quRcB/pzwx/1Du4EpgPaeNII/hhdh2YqBY8LqZ4bT62Ig
NC5p4IAbHsLWYYGCHBoGAEI691VLtaXUUcU+cJ/Jo8gQp2dgfsTnWvrIW3iXnaSkjaldazDnR6c6
LInJrPjB0HxqHXpYTmog9Ef4WRerZUY9leYvJFc9BsEek9BdrqSXdoeh2XmwL6M1wK9GTMeFTsry
VgQedQa17AsK308wpNaql6TIQnIRkmf6/wiQPt9UfFou5o+3JFiCKGTwL0ouCh85qJnubwym9Eu2
5FLr0VL1RQ6CNmYblV6klB9g+UXfKn0bukkcjXZuzZPpKVucmtqXeMRh1oMEpdjspXSjOfU/gcND
Hkp0nS4l1SQ3I2NapkBozrUxONbeuTUFqI3apj693jsWgyHAb6yH90yNQdQcM6Pp31nV+eDmdHJK
AWA/zwzXdLKcsF6/+grPgr21EvEs9+flqNE1cLRmA0DVE5eWYwk0vhTXDfzkQmN3XgPzN2v+Crmb
Xw4a5YyUjRuAQK5/WcNeueg33c6wvySkTSp2+cKze3FOHPjLBoT1USaYBEywf4b6FrxImkVLFoWe
GR/8pEdg9yTx+IAeGCU//YBE+P7+UFTYq0op1IpW9nqBvcSteKXiAIb4QqCXYnBNwJzRD9ASQyMx
onx+jJVUlTC7dZj9Z0JbfmFXRv+Qp5ReZaTUHO+p7g5p+g2o4eRTW7FbgvTuHRrmDIT97qRqwCyz
nCpZnxoE+xXaIqiQZGjmDaVykyUc4/qEjXIcggPR5bB3nGDkrA3cmT/7xWoSR3b99vCXe+/6UMZz
WlKuSSGakRscn5TA/gGxxvnQ6ksupQcbZlj0RAI3+GvLtaBVBR2cMeCtDT3j9WJ5vCHxt2A3NzdU
swccYCiO+Bdfz3WRZ8rH3gy/duqhSmfYfzhBphGDkUxXrjGdw8g8cWMLNhpEErPLthMd0VktiBAm
wKbL8gfKD5g/v8nZhGxZFjNGt8zw8yd6/qRm7wINDlXwQo1C8omZ9lLMDc2lZlXbjU4yB5VnCVyS
y7ZRcEEC7qbINH2CvVjyP6Mja0EhTfesbc0QSN8EZZXEkMTfART4tG4TDG9fzx6gUog9J5vFZ1y0
VOovvylS6vfiDhugtZaifwtH1V7rNNL8D9dCg9+N+HIcWnHPuWrZ2mQGofLK8RXgef9SiQzwzdp7
ENkMz4OJ/MJJG5OvDyFUjorUZV7LSX2yh6vayLkozesmqkla+sKdriX5QpeR2xQlJxS04sWodkdJ
mFVEiyzwrpGxEnR+Cbj1fnxi0lmoEeiV2kGNPtUzbzNhcS+B0MV6ee8l8YZNT17moWzx41O5JfO+
hFBrgpD2X2yDTE1VEHkhn87KRCIOTIYMDK2tj7PzcxQvNzaB304Rw7V4QhJjvNezUzWfHcsrpRC1
her/whqtztcOEaxS3N8GAEaC9LgjXKqmTfo4p8pNjXL+Hc5MUZgQ/loiiYTR1j9/JmriEeDhAAuf
mhjj41p20XsPSY6aUph4JkPlcxx+rCtN1Cf+OpwAOnrpIA8HtXEpWpIh6MDWXLzO6wr+MvUsl6p4
+EOuMlAK16D/fjC0HGR3x0VY7l+M4gNxQxoiWUJ+yWD4v3dBauQKcZuG7YqrZOn/09lCmNBi3H13
MYKbd5pakRMw2KdHaRjtVEyYYlSPedOJqKHVdLRMzeHwaxfJdLjzx/u9mzlS0HSe7kjDUsIbpxly
7sK95QkzjvIkpKArkiuMIfkce0fbBYSx7TV3Gr2UxLXIxGapn+3lIYtmQpjDnnKunulBFxY/9xWE
Wya+Q9pygkBkdGcdE7SYC+koYVsRJ7jB11PhkVWglj2ZWSgBqLzmJzbjIymqEX8C6AQpfAYgUcc+
5B2mKphgHxsvfPfkk1hC5gV0T/miylAp8HPWDqtW76OPJzEl5I1pmw3GiR3UPH77WRp7KKPKca5Q
ggK9t3WLhyOX2D8Ff8cWZLZuqcyj6YWjPhfhbX0R/wfBkxMSlM0ZUM0MGvSUi1siS0R/bQ1ar1tL
3GJlB7M8rKWNREyBCxgoSEnLiRBR7yyPwWtnqJNo682PjPBLTfQMP6uJAx6ibeex1p3HGAIUcdQC
WitbHgyzraXQsJ18KKkqV0xDyR8YNMtajUHq9LVPWlIMaSrE6lW3RqpBe4Ey4T+v2VYK62DYzUZP
EXNBzanEuneCg/l39rqBiTA9w1pKRI/k1XIkYc9YJJu9k8K3JOyDucJxizHjehRzUQ+tUV63uRFU
o/03mzzFKjSsDYRfL/Y1Vuq4fa9qC6V0j461oc4R2PNqLYt0x7eXpQ1PdZITnUbxaZzBwbT6n9sE
FfngZl7AR7lcBmDlvLZ45hpNWw2qQ2d0V8ZqrYLycu1maIARGN+QgzXHXdWUlZDhGKBiaBM8BLgA
OtjEVUCp4lvmr+LYEeAQYw3rH0tLvWUCiHpH/G0oqWvukd1kBvez0GxHwz9rj2p8kgYga4QCj9jU
NAGP+BYlFAfM6e3cNKX+jtV2kdJAxELJ4M3xkHslOFkTyJiy3i2TTsM9HEe6vgsUrcM5g7Uw5E3R
XrcSnp3Tpd2E7AkG4pZGyhjGtJp7it6vYZGycc0AomDKl8DLjOAJ3bOly7VngoI9sDhbK0lWgmgF
ap95ChqEjYvGgd+P5/WtDWugEFXT6WjSc/QACzvs+i0Jh60ITmY437qm0OEKEtXzdaPMb+aD6lXM
byu+R5i8JiSlNwgxvE9hObXb6nNQb3Iqr+U2Bk1yGnHk54/AeWkMganfVLNz0hfu1ogEjefwoCkE
RyfQkKbjYqY2JapK9MbettfzAegrZhgsPE5p8luNWy1JJpSArU/5kXVLXqCvomfITiz4xyAJxojT
Nf7/Jp27EbNy5Kdazvx7ZjvnKhmh9SpbifgOaljDMR3X4IdVP+6RMqNHseYqaiZFVH+TlQo5oVaf
AnFPN7qRsSnd/9Aad2GYyaAnP698hLemKytuKxkhLOQOuyBgP67eO1+7t3IJfWphLQ9rf4+ifGGW
NtmQUyqDpQwONhhfcc5YH2lza/dUObq4Ezp2D3cJ593tEMPTV/sljt8mv1T4JJW1QSDgX4ewVMsu
KL0dEGsdhq0jsIviRNIk8moW8yPB2MW6lVL0ec4l7+h1zge9G9upkJ8hOKHujzKKBc1HMHH3DgtF
3DFEH1DhM4Cq6Xqk1AH/+SAghFfrYGyeUIkf9Uqtp14rbNR/BmoninboOTiUG/KbqZXshuPlNwg/
LO1Gnu5VhSNEbQreL0Sd6uSPPxi3MUcEnj0ZQt4M/TcSS4k6FkX2L39tolBeVjgBr0e8hZtHYiPr
jM84GtWwL7dYiByW8S4JVurBrb95X0bc+YoJ3ZC84JeFkpbDt9iDsGrqaa+IpihKTOdYwKp/FxPN
T2fB4W4WWWuIAVLLNR3k4DFO2TXUqtt5bDpmyHZoBYuzomj7rFkII1kn6m1Q0kqty2UCs3HSx89p
QebuolvJjVP6AcrYspqQkpjKfAM0omLgcuvILArHWvZ3kmClMz/JR7knSFQVpBIBPKo4xFoQkIZh
jC1nStP2gqnAEUsC98atUF6j3f9fCrCEDXm4wCVB4UjLzQsbflV8a4ED64hkcWvprEKX2cW8LZn0
X8Dpv1B+d7fHLPAcl8zor4YS3yQ/jeeEQHNUJ0nu9RplCVovcdvnShpTfs4xivHix2yOqSvhgwgP
AVEmqF8zkeLhGisQtChw9ZPbhl71fy1nw+boAAbo8WMkocfYwKZZWHk+Z3KZHcjwzvGAt+NI42RH
QFRqvuLlQ4lK/7HLATI9OhB3L46/eW0rIbZC3rlRjFKsZ4uQpQjCNegQWV+Pwn/jiAtAOSNHy8wr
kgaJT8YqLeOF9HWTBhsy1d8b/vyDVlvnls6WFa9ugYvwQdd4QgiPilEyEM2xOKLFgrPqUtL3hThs
nX37Q0R7w8BV6t/iR1dJAL3SJSsZUJ/oQm6fiywVreUH9I18IJvXO+rlpmD5cKMqwRXyCNNY4/ON
8KTztmOkU962iLm6v7dtnth8fVjJhc9KkFuX8/DrcTK9wZoz5a7QV487ibNsBNq3hfeEupg7hPHg
ShFdO1TjzI85h7Ic2YyQ9HgN1lvRHzc064Xyz9O6n+k8Q0QJgoh8xT89m/KqQMp8ks243V/x2TfU
z8KNdByXDy9rjqTCsoCherE2IuysMPWrc3580EP3TBjcUmjcu3I5FV0UO8r0NgW4xHs69K3ejU+l
vFND3vCC5dPdbAa3Hx8ZTWxsAsBolp6Sj06VPCjN7erANZTfwXF+ebqartbmE3eH5jgUGbiVov7h
HYklKF6LXXTtag6VLud6sZr/yLS2qYAaIgduuA==
`protect end_protected
