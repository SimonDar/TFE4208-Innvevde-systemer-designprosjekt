��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U@W~z,r#��$��ٙ�����8�I�u������^>:��JVҌ+�w��1�N�]�v�[`B-O���[nT�<���v��QR�Wf�R`�d�@M	�'�ؾ�����tr�%�^b��f<�����}�+����m ��!>%�	� � ���A-*�xke#ن�f�}��h�b$��~������L��!���M&J���da��/ec2�j�	�s>�B}܎g�3�j�t���q�[�~���uOa��6Ca(`��H7g��]����]�����5K�bS��2���¹6�Β���Kͮc�4 ��WE? b����28Ļ�:bW�����ξ��,����
���<���X
������JK�F�`g%i�����^iC��n��D˸�\jҿr ��%B(}��Q����ʼ��r||���ȇn�!�I�v�?�N@>�ME�Q��<��/��Y���6�4��`�'���1�.L�+ض�[��+�X����-n�䏠q�j1��Wbp3RWG�������JJxa���;.��=�H�4��ܺ��j�	��Vy �*'��q@�����s��~���O�!�n������MӞ��h&y/l/��u/2�L y�`*�Z&w�c�q���&��q��u!V�
b��,1=�N2ʦ'$��S��8���d�t���W+g�	D�m��� ��'�ȠPp���7X�Yv_ߘ��xO���Ã�b��@���	��3I%0���V��d��$&3o���n@��}�2�7<��r�K-r�L�w3Mq�V�����X�BR乲������Kc��Ԩy
�̐V��35��3���� S�6�ga�&��H�etQ?�z��M��,<�!5:IZm��a��4�Cd��yRQ�zH���i�8]�`G�~Xb���z�v}9S�r;��\�����4�@��?�|wG(fR�&���&{9(+�dka]�"6�	D3�iB�.6	*^%�bZ$�Λ������o�� ��|�g���e/���~�.k`�)w%�$'Ec�$�2����hFx�X��*S�Q���ƌo�D���:3��t#��X�æ��q,)�����}��
�c�����H#h��{��P:����H{��r65���:	E��r'�Q)��qy �yh���gg�V#Z�|�n�|g������-��`�49���V��R��2YgH�hlM�A��O@;��[2�p�3�)� oP֕��4���\hh�/ǳI�_ݚ�!��{�Ćg��0k�9⡊��}!��GQf�� 5����oPv�*\m��P�c��w�Uż}]gqb:��g�0EL�x�u�����<���7���Z�}�O��a��ez�\A�c;h��j�D���E�@/q�Y	�S;P%� {�g&e���R1��2j�!e���\60G��֦*�@L<x��L��P/���R�p�,O��}~L駿���.WLV}$�LA�o�ߊ���vM�8��I���J�x=�](x����~��k�٦�C.9�^�OX�2����R��)��H�oI �� �&$Gp�ª]��:QK�k��c�D;�;�3�|���l�F�6Ԅ�}�2<f�}d�~^}�0Pp�l�k�:�6_Ww�V�T�����ۍ�ɐh���J�cg�T���md�?+��l|��<���NcG�i�ԍ=ާ��Is��?}�$�ں�\�gY���'t!��r;����&��
˄����w�lek9ӌүsx��u��*�D9��y$�@i�xi�]��!掠��vw����bqq)Ocݴ�M�_O��<�1*�JϿɮ�Ʂ�N���Fj���P9�L��z}��F�#�Z�� {$��i��1!��\�&CW������X���a.���pGpJ��ϐ�c��n�x��҅[��{�����7�����U�B�ݯR��d��N5�D�v��W/�|z�����upK9��!��G�Zq���V��R���2X��l�o���1�kR�HY�f?����9���J�Sd��ʃ]R�����la@���2�a(�f���('�L����|�tB��J����w&!Ʉ1��Z�>�*W�5f�[�?�5An`�"d�BHy2��
� �'u��h�\[�z�r\a�Z����fɹ4!� �u����h�F�=-([�V�IJoέ0-6=i�f_�B=��d�K
[<��G���bW�Zx#8����N�/�>�[=�����Z(o�d�\yڣ��+4��w���s��C��'�s��~
W�3�7�-���<�}ֹ��Ӝ�a>T��&�\�'���h6��n�;g4[1���[HI�M��U9����q-��A��3����k0V�����E�"��[����M�RK������x\r|lU�G��L�~z'�s�XͿ���ݥ�	��6)��8N_X��JS�ƺm�MSs.ȡ��#�(9�;�i
�F���|j�8>;]����fD8[�����P$�zL$r*vkR��i���
�
��W��m�� �56�<���
x��쨹������rl&�Ɇ���A���e���4�������'/�0 T�Km�
a�b�a�S	Z���x%g�%��enO#�����i�D[��]Gf5�H2��ì>n*��^@�����3SǎS��Zif)�ٻ]�x��_�	:�` �C��^U)��&�U��۞�*��=r��0)�&)��y�ؔ��]�k�8���x�[���v�p2�g��\�^#D�ۢ�ú����C?�:�:������.����3\���Ap�/�7 �7z&G��8�� �?�j.$ܕ3e���GIS��hqP��3+B933�����b�C�۸k�ʼ����C��I�a|�_�SB_#8��|z~��,��a��Y���_�}���j���R�(�	�)R ���X�L�X&E����jt��]�(�/(�G�F�Q�J��lh¡��̖��TU�?�=������q#�=�����5��X�CV��|����p�����pfݼ���:bp��I��S"��Y	��7����td��ڎax��XG�b�!/������ك�r���p��lu���S��T��&��;�X��C� >�b�|�jw�9 Y� ;E zn�Q��V�E��-B?�M����	5�)����c��0�*w��#�<�cU�2sђe˕sk�&��F�����+T��t�gNɡ�;���n@9:�7��(+�<�B�\#-�;0�(M�*��>	�U�2�n���1[���#*�����������x��0����I��2ER�Z���ns���%b�����FL�h���60�$\-3KrP�Q��3 �(⦐C�8a������Ǵ|����R`J�y�V]��b�t�� ''�*�v�;���1P�㸥fMA�yi�0�P.�0BƊ1���7�wo+B#Ȼ�7����抽�,�h���C͏���u?�Uӯ�/�6���l7Z��@M�TO�x��������p���"�������cN>zg��u5��V��!�nu��鴯pHw6�*�wIi�z�v��ۻ����^�Je��'o��-�֋�nC�E��:+Id�Y�C��dwr�k��˾�ڥ�����bۛҴ�%λ�Cg��eK��ǘ���V�v:4��Tk�e�g��oU�HH��0��;�v�NE����;&	���y߶�%�34�i@�?~��b����T�o��<�sLV��[���]J�]fy07�e��cc���`�]7�Yo��������X���%+O��YYQ�MM�tA�⏌o@�]ؕ͘vY��\���Mwg�[�:Yl����h�8ψn�g~��>���p:=�8���ܒk��P���u/7l��旺�m�W3����X�O�����sT-j�H�ר/OK��*|�*[�!�<�v�0�s���ԅ1'*����'SE�=�߸(�Ԫ��B���`�R��ޣOӴ���l��	;:��w������,(���rR5����*/~���Ҝ{S���-6V�G����z\��Q V�8��S��$rN����G�dR{f���ηpL-�ұ��U_���%�R�Jk���g��b�r��'u��6
�³�����YM��&�{c��ѵ�]�]f���ڏ[���V�M��)�B�S�o��u���:
i2��2@R��x�0�n'��GY��t�`Iͭ>�O=C8� K,Daܾ��	�n����E�+�g������V׃G����/�A�� ]�*Bt����=u,Ȃ3�6���{���j����W):!\Ԃ��>�X`�9k"W><��s_��ʰa��{))m�x�Ȥ���'?��޷#RSurk�c��f@c��WY ���r����_��z�ϒ��N��R��<�	��=SG��ٛ�U���]Ē�B&gW?�4�� �6h����a������K�9,�"�w`~]�>Kpj�A�C�C'W�L��?�����A12����?܋.x@]��6�!u�U�㊳�ϱ@�o�;��n���b��Ҡ�hR���g���O���z탛U?�ۦ~� ׆|ߘ
��T{�}�AE8�^4.�Itgp�j�R����%��nQ���_/�<�*��d��Lu��g�sP�;�F,�R|�BH��fr��۫fV����o�� ~���![����t��]W{�n�� "#`����)�@�d����l(*~1�zJ��H1��S5�(w��e~��w���3�������v@~w�3[ԣ��I����L �I�r?*9�R����x�2?��]�����z��?x6P�Z�$uG�(��籈wx*�-]�D�&d�����vM�$��g�\`�G'x��I:�`7��M��Aj���m�"(�S�>�6h�W��=|�I��JD�8�?W*�����BpV1�_O�X�(�y7���nl<E�m�|�ߞ�V1߀b��<,��
��r�����X�ͣ �f���	+���Z[!CϠ$NOWo#4Û���H��8�+��=����ɴk�� �I�zYC�ܣ\WT<:�!?UIpv�*Uf�m�����[� �㇡2�F+�(N�0|�>�u4�'�}�x_� �L�-f��1�������۫뫛��)����R��t��I��~�{(�,t;>�m��fN.�cn�b},=p/:=�h��'��,��� �Yq&d�!�����06[bp�	��g�Mv ,� �k9����%�H<S̿T����y��v��FޱP(�;�����S���hbX�Օ>�mzK�'�N�Q��gs��H ��}ĭ�i��VI<1�(|%/T؃B*�h,�c�<�+����\������.�g������02"�S"1j��xqS'�-Ȃ?�b]�h'Hw0,\n7��I�H�{g@ �Q���v�)�#8s1�!���$�t�_+s>��Ǣ���&�}h,mK7Uv&��陯�-��[��nA1�I@I*\Ɍ���j2P�M�h���I�}13�� 8�����a�a������\��	(�d:>�GOÎ�����>r�ܐ�������_zپ�b�f�'��Y�ރ5��;�g��Èר��7$f��1����y�(�����#L_*=E�ĵ�9J*R��C���-�q���X���☫��>^�~m����{�* S7�f���R`Kߤ�ճ0�P�Nʱ���	�����_��ח$��H)�y�nV{p6��K��mZ)n�hA������ꇨLui�\��z[b���$�Y����`0��� ��5�5���v)8�!ȼcÆql���/�# UDVb`�W���u���T�4Vah�7�q:X3�Y�YHV+�-#x��3yIH<y�A����}F��ʛ�{y��<� #�b�)/�}DiɹB �8�2�g���!j��P��n�~/�s���E���X�)�dn���h
��������\��|��;�u�j����e2ܡ.khA�'�����Gd�k!��2[L-�!Ѵ�Y�<i1�:RlRGGi��R�-ZW�����~��s`;h�X��x��!@���%\#����:F��F��(j����^bZU� x�ѻg�<1��;��K�|�+���zZ��m����Z�F��Yw�*�	�`�M���o Pnn�Ec�P�}��D�#3��r�_����a��X�F��|��;RV�D�/J���?k#F�8�2��xzu)�\>`�t17��z7�w���k��` +�(���Bv����������b�H1�������M�I����M1C�hj��W �"  6l�0���+��WJ�u.h�a���Ŏ����5<��3�/ \���@�):B5�w��ƾ&�
٩������#��tH��s>y�{T�<��SH($y�s�����kh6#&�BA��L���8]�9���H=.�J-����hX.]l4t�O��"���k$4�{�c�R��埥A�u��G�s�H�|��r����*�ak�#�#ɬ�k����pў�y���`��2���͂G���՘�VW�;BU��X9nS���N�o��*��i�7���'z{b��^�B@ a�+L` �U++��������������W��άhfze�Fe�"�g�W���؜`eی��q���d=����7���kXo͙yH"Z�^���A�X��~��� ���>>7-H�Q],;"¦��d������Ȣ_���Wn��+��!��m����Nƴ�CO�!1�j�'�Q ���"W'���|?ɹ�ł�f$i�5g5G[>t$@��.�r�@[�n���������p��Z��zM�󓊔�_ i��K!{��<+��t�/g��E�4S����X�b>�ޡ@����h�76׶�R(e{o�Yl��>n��h���d��_s䗕� �Ŷ�Q:��|�aS�
��V?G�j�v�:&�b�U6����2��a2-���@�{���χcc��,�z!Z]�1�aN��)��e�	�a���Kxi�-8�»���{>S�Eh�lV�P ���ϭPo�#ua9{Q ��;L|����i�mLg:�zg�WS)�qiC9%�C\nf��/x-)O���G�#�T�p�	�E7�X�)�|��<PCk<4�3;R��eA�bh�I��qUرX�޾�F#���t�������`�I���m݅/fC.��a�ܚ/u[�'�"����ؖY�!�. �Xv���$������*qd����C����_��hO�~�W;pR#vX�S��/"�"W�/oV#�P!|=�,�
�r��5k�nu�c���0�i��'S���z@���+��F���uq_]b�kz���b�����8shG�)>�̥=��%��1�18�syw�JIy�9�f(�l��3Buِ.�һ]E�+QhQ�Ȃ�3��I�uᙓګ�Υc�Yֿ�pM_�j�i$��M;/��n�*2�g~i�.��fW���F�rc�� ��5sy�^!{T������p�J�'"��T�����O�^V�`}Y�P�?|20ԅr�u���?�)!�y���#��Zw�+�M���>�����)b�kH�K��r00EI6 	OXZLZW�e���*��Pr�q	���DjÑ#i�.��D�ϋ��ͱ{8��&�ym�!����B!\�W�c#��j�`����g%��<"��M��nt%�J�v:�Ӑ�v��aר��GG&Uo���1u� ߺ�(���7��p���[M��޸�TGz���6ư\��۟�/a	1kf�h���~�<�����.v�ոxh}�LP�iʜ_�����������^y5o��<X�A�Pq,#p���⎰�?]`O?#zP��RT �jbS
�����ߔ�p��2]"I����˥Ye=��N睯�O�RL�	3-Y!�7��c��W�Ϋ \{vG�y���B�:�����e��]8��tj�!�I(��v��=)�]��R�C�n���b�L�0[��POO{�'�sڐEB��d�(n+��`:�I�S)��^��Jly����-���#E�3=�@0{p���_���}j9P��@O���4"S8�����{��ew���l:Cv�
P	��.�su�cPĻX/l�g�]����)	���̻��r-~�rQ���i_�Ү�,�D��&�Si��~Y$��$��ğ���H�ח��.�c+'��Or��k����M�L:���7�+H������)�V����7��Q� �#%��B�;�� Ux�s��; ���¬FX���z�[�j�Ïg͢��%^�#�9��nߏ(�v(j���'��
fw
��6�bZ:[\0�c��@RK0�Z�� �8c;�P�A����i��6k@̸/�T�c1>F�b"�[����Q��S�:<��JV��]c{~�<vtǡ1P��s�	G�Z&t�uP�%o��K^񺜵��a�W�蔒S�F�{�����m2ڝ��vxLRe`�O�OL�����[�»f>Bqs˅��h���������q*X����1FPc�͜p�lx܅2*(��i#Y�*���_����{����6��3�
��Ο��D������f��ǣ� AX���I�Z9��xƠ�]���`��Ԓ{����JH��o��d1��j�� �L_�F;^�}���P�<^䭻�����,/���Dg�hQ��~Gai.�!����
�w�~�V��>���9Y�}��J~��c��Ơyq�)��)���9�{Q�P�<Fy34�;�06�jЃ�8Tw�y��*���P���}�J$�7�Ņ}��t��}s3g!KI�୓��n������֍6��1���Ȳ�7���tI�.ώ�DP4��[Me_UԖX�Cq&rE�̍MU�ň� ����g�.��n���[{��>���3{��������*�ܰ0���ď��eO�os`�D�M�Ďz�½R�;��!PF�����^|�1]�t�Zt
�k�ο'���OCZ�4�ʦ������~zE�C��pF<$��\�)?�Es���/NШ��*,�Lvf3�gߎ+�Y˴2�r}��	S�y}Q9 �Y ���2�f�h��e��KEhk���Y�T����rO�0G������	�~��kH�~�k�s�F-��"w���������n��ͳ1�%����j�����V��WH�X.4�t&�����X���]GK�!A$��� ��T�ᡄH<g�L�w�R[�T����5>I�CR����?>�74t�l�<��o�p4=ڶ�'��ߧ�c�q8��G�q0��$濰�";�`az�����y��^f=XXYq21��%"��=���*)����
�7�2ꖍͭ��F�bVJ�^��\8mn{jͲEmo�F���{5��hu#s�MhоcF�q��Dn����J���T�<��Ś:����z[�4��Q���Z����0� ^�F߯>@��{o��M�A����=Q|Ol xV�O�(�^�9���ն{B=_G��k�>��fϯk����HL����j���y�[��.�fv���zq�{V�EyC�k��<ٜ�N4�x���W�DiF,7͚
Q�D�j�|��-� @� ͮ��Xٖ�'�>�泫ց���\=�Ԓɳ)q|����W<�|O�ʜ��+��ݡ)��naK����t� �%���"���4������sc�Dkx����U�������TzK;��x��Gj�OrM-I���A�] ��mi5u���o�_��k�^��ʁ���Kq���X>!����`a)3;>V�0ƨw���{ ���E�]�h�+I5��]�Xص�r�&N��\�&Km��x�x�跦�7TTw���s!Mdf�-�g!B'��a�-��r�m�9�!³�z��2��A]��d=�������&$�_�.�ut�����E�^;�$X �̞��j��2�W��^�9]dQ`�T	�K�HR�GSǷ s�-��{�.� q�{��ԲV�3��"g��$�05`4kq��SVdm������2��
m�x�=�d��'�#��b��SN��g֫:�9i�c�{�zPY-��i���54���" �ֻ-��_	K���؝@0a=rߔ �KoKL{���Z�h@���(VZ��(�:#���L�V4^J�;B��U��A5��-?��� �����|�Gh�� ��:�GC+�G���7sn�C����KhL8V&��\R�S�3۹4�i�MoA�#՝�g�u8��ږ԰wi�d���gO��� 2�nV�d��2������໡oqJ��;�}�g�Q�6P�V��>�B��l����V��7�w������!Lv�M�VLFs���^�k�;p�ʵ��3%��U�T��e_���>��޿�d�ʭ��������[C;-���$�-�B�íc͛\�^�w�̩̽�Tl��f,��[r]����aض�C����q,3�3t�����1�m���ݦ|�5,�d�"�
r��={�0?LT�	�FW���;�3 s�|�xTV�;C7��e��c��bN�����?������K�5���Az�:���S��%T��.3�8��ȿ�̋؃����qUs[� �W=�"���
E�"��z.��e�j*��J��)�eO�|�z�М�{�ٸE��6H��J�ihO_���(q�#T�_�� ����M�$*���ЇC?,7"�Y����+��=�UK$;���I_�F?���2�*���˯d�*cEs��S��"DAZ�����HGI�2F6f��Ϫ ǭ��v@�zم٦@�+�9��u-�n&�p=R������K4t�(�$��m1�z;-Ld���L��e�c[&�Ӕ^Z�Ck���I�ۦ��_4?p�Ҫ�.���J"$.hxyġ/ܻ@�n�u�X��]W��Y�}�oyCt[�M&�[ŭ��Ԓ���*2*)��hb��!�(��J/�Ҥ3�m����\{`�d ��aJ�qM�B�*N+�	k���E��y�и�5��?�+��h��CJ��HLK�&zf�A��J4�� �[�#B۩{�oz�01=�j�����C���Y��m[�<=��H��gF5S���+F(�s��e�42�#�[5�ֿ75�D�]a'򀉳���O+c����7镵�Qe�Z��0��$N�ĳ�sQ����U�bB������'�·��.~A;K�0�^���QI�ܴ��mW`����@���6J��c��Ū*�lB9}�4�?5!���MU�O6AF~����M� ׇ�KP.'����F��ǫ�Dl��� ��C!,�$�¹�z��	q��M�IªV��}J΍���=
�]�ixW�E�r��v��4(�t�ĻO02�A�Z��˭�ۣ,n�z�5g&{����vGlxg`�ւV�#� p`,U.���`�-�ا3��ʠܰ61y�])A�޷�;�n��V Y�2��u�
�t�UF�a�v\մ���f!I�y�B�c�]v�t��рgB�{Μ\W3d���&PVp*u��[y�ZX|3R�1H��8wWT�Ii�}�'4P�}�����jQ*|�����n5G�
���*��L1�:��;]3��̒�*|�������>]�"}�}�J�K:�!��`��?�A�{�G�"�{n0U�!��F}��l�zy��g���K)���B�蛧�$r�o/��@��ef/�3�`W<���G���BN����$ѷ5Ea�p5�S�[V���,.|�S[���g�͠�!}[��K�ls�љ����f��X�]�2�*eԚ���
F�'R�W��T0ߞ|��j�P|m�Fo�������'�U��~r��g�P3
�*������]ǏWLg�e�i$��G��f󭋪עG����O\�\\��ǁ�'�W�^���i�"K��qxٮ,&���s��b�姖'�2�C㭖��q�]�,%C��$Y��34��y�.��7ۧ���q��|M0��_;�rNm�Zq�2��cO��<g����B(��[�v�z��
o������]��' ��6��n#H�ϳ��*|C���L�2�%�p��NZ�GC6s���S�6 ��y��Z�6!T��@�3��p����]DK2�o����S�狥��<�Z}]eɪ�H�Y��-g|��0�<��O�#;���U �������A���\牎~4n..l�+�B݊�$��p����i>�]��A�� ���'%<S�]u��❶����e_tg���:�F����>��2'>u];�7�ƣ�ퟚ wH��e����M6H�x��s�^=�eD�{ʲW��u���%O��
�c�#ɕ�tVZ;��=����F��R�@���9]�KD�ZT�����kJu�r��@5�}]�g�L�9:^��^���-W�
UB�-���;�"�jr��ķ�_ݨ����A{q9�Y��T�j���NYi�j�'�p��<�Ϡ�K���H4|�^3i� ���󶞞e���  Sv���u�O{*��@��V$�Z��V"j8�h Z�+����p6�ȟ;b�$��4��|$�5����<�+���v��`�+ޠ\Q]䢉��y��X5ӁU�'��g��CHAy|xW �NKA���S#�KFf���3�$���C��g�%�8r�;�'��L0[L�1c��ހ���S@#��w�
LLX��%�Vt+���Q�r9��}U9��G%�ԫh����M�#x��ZY�*�Sek�}𓖠�
q]-_ �`G�2ܛ�Dܜ������ZLo�zc��X����,H��:���M����i�2���š��j�^�0��@�}6�J�LY�p���u>�H�U� R�?�6k��t����Z�U����E�m�~� !\S���)+\4+fW�sT 1-y�i�\:1� �J%POp꘾��'�z;}�!fn�ݙ�MT��%JGK��ɓ@"Oӊג���<�~|���n�もp�W���{i�Ѭ��z+�ݺ6��b<f)z�UV,� �X�����% ��z
�(o̚���)k}�!j�\�m4[5X,FS,b�U��?�7���`y�0hĹˑ����A����Mh��p�oGD�V���`��w._�$|Ld��9*ys>X���2ȯl؅���d��`>��VB����/Ѿ�e,'������P���,x��6���2+� Z��9�	�qc`ߡ��هxr�8U��]�&3�ml�i]A���\��O���\b���vp;$vTMҺ�#��D0���˩Ĥ���z�P5s�&lc#���[�A��Xw��z'�����4A�!�Y f����ﵔ{�Z�U�WJEc ���H!�y�>�s��T�,��.�!�N��~�>g�=퓤�?S�X�@���B�%���������������g�t�}u�x���ޙ���O�t�m��� ��MlH]%��㽻����G���9 �E��ԙ����y�ЇAV�V+�,��
��~��Ѝ���?-����]kV"��͜d�糜�^�jH��K���W���w? 4�ލ�o�8�m:D5�\��mg�Bmz	v?�w/qvG(9�rIb�������Al׷�YA�V["�ľ(^�U{�
��4:R����[�Z��bA�Բ}F���^�=��$�����j�W���/P�I�A�{q_K��Ϙ����l=$&�!�kP+�-hŽP��F:�5Ɍ�.7��F��æ�#U�����&`�ɉg�oU�aW`�s�5Nn͂@��]w�����H�����W+�-W�VE{��C,M3y6�[�.(�Y3��4����@a�O����+T,�L*�|8�����*n3![�;����I�1�I��� �cc�Ū6�ڔ<|��z��J�g���M-F�p�/��V����q�<���4R��C$�U��D��攨}>q�֍5��슡8�vS3��ܝ�}�젹�%ffE[�%�e��xpaZ�E�K�_���.8£{��k5���ϔט*�N�f]���A�fƕ�q��P� �P r:|��%	�����4!����I�Q��-o+�����*�<�;ƴҢɐN���\�sR�M�2�������aq�t��Ȁ�_X���ԁc��bz��ث�х���N��%��Z����̔P���Ǐ ���|������),�g����PJ��L=�G�T�"B$.%͙�5GB�9o���j�?��y��l꿶��~��n�7� �l����]܃����EP��%R	f��6nh"D�EA��K\��a5MK��[��c@0v�38v�^7��}�G�R��%��䌜��b�/�>N�5�� ̹�[/���Β��^�r���6��럡P	�baO�O˦�_�W]zc'�"�-��'�A��D�ԭk�й*%#�S��E�<K�=�S��C�N�� ֑�}��Kɮn=�z6����0l������f��-,��{��-s�̇\;���p�?K�ެ��2)�⿇(E�Ē|��і%U��"�3ܼ���v�R��\�[N2����x�K�:�730ޛ��R�K�O@���5x�Y����K�H��H��!��Yɹ��Ӊ��A��X[�j��W
34�.)��D�Da3���v"A�98W�u���L��w�;��RAƶ��᠀~~s�r��׺y?ޅ�ң��9���g����U�#�u�O������=����
��:�]դ�5̣\�`�=��>�X�,��[���̺cqFG\ʞ`6�$�C�A,���`��5�ig� ���e�O� /���7~���R*���|�t�|��;qP�1l'�t�M�$)m����shP���u}��ԕ,.qR	˨\��P�t���WH)�n�`n��ќp���޲'
�'av���tG��/b�𮁴��ח<�`��=�r�����E�0�.�1U��q֨��fIc�4{�j��$�x?tOؼ^B�h�����i����M���E����	k�Ew�P���M�,�ϲ(����/j���8P��J����6g`��Fg�?�"��8)�^��2��v4�1_5����F
C����MA-#���y�T�;	8���Ⱦ�`O���bE�4M�~e�r���}�H�O������Z�YT�2�2�w1\8�`�=��.|���o�@�2���q������$_�gZ�(xq�U~���C>���<#���2��K\U�{�}|�QF�:�)�����݋^E��&��Xo����ф��+�)��?6W���;�0��2�
B���ޔ�*}���{Xh��\��q��g��V�=�\��7�*����r5G��h��k:]���BzI���<�� ^��
7�Í�1�q��薶�.�Oy����^��L
����#��Y���9p�@'^���YSu�M���D��w-m��vEI3�ZI g��?3@`��@�����g6�ef�#!Yx��4f�U#����gƲB�/St�?�
q���w��"�Ԓ���B@���38��Z�+X�~chD�G�J���f� a�D�����'��jw3d����#�#�3�J��m��7C62�[���9?m�t��ݻUtL7/:�>�O��O�\��.˃xzW�����R�zj4�#�ӧv-H����e�Ȗ�B9��g�l�G��-��!���,t7cȎ���\��ؗ������r(��\�a��_$߻*�$Q�:<Ip����B0�"�����"O������E�NX�-�N5#��N0�k��!x��jH>�n���0B5�����ԧ/�6��hU��� B�D.����C�*��#�}�bW�`$ȱ��_͈�5���\$��ۖQ��e[[��e����d��������Ä�8ȹ`iU�������sY��qNg]�r�_"�5�6XV+�>�u�;`h����/憟޲c�#���"�h���
��ؐ�Y����7���l������#!���ㄹ�6<C��d����	@8V�{<��J��L���j��C�o��Wu��IE�[�\8�m�lM�x�����W7��R=�?�ڧl���^�:}I��<�|t��b�d�(6��`���L��z���|:������5]�d5��֝��Rvba�dG���a��<��F�Gv��Bۉ A^K�.�nBgC2��9� OWUI��x�8	HNm�^n)І�ιv�GWZe��_�V߯�)֜�Kh� �O�!�O��Mg9�EV�1�a<Z�K۞>D�D����h<K�1��܍�ƴ�1Avii���uz�;z�vf��Q9G��sJ��)�{��
;�ORY�{�X�y���JҷV�E	k@frZ��k�W�V�%�׍��/�����є��I�S1��x���h�!dk��A(1����^{^���B�>%���~��n�ڬ{A�rѭ��sB��Am��'bCf�5D�2&a�G�q�'���A`@���Qˑ�g0�f�M��?��V�"g?�_�m��ȸ�B�& �Hq
����o|^��µդb�T����u�ݨl�W��<K�ʪM�Z'0=�d�{J��#knT�:N�I�3T�U�I��:{�c�s@$��f��jfTw�r9
'�'URN�����������N:�®�d���ܡ�J�~�h4�����״{���<��gL�yښ�f+LisZS�u4�ba�g�̣x�$♜t�^alg�%'ZYaʈ	ŵ�}���-�+�"�B�L�\�����]-we�	�>��bwp�%\����� ��_ⰷ6���p���v���
�BG��=4���[{�b�sj���$ ��xe���bs�����1�'N�t}(��4a!��	�b ��F��W(�PH]������UI�i�ҊB��q#����Zt�q�G�l��X�PU��:r�#߹��C:>�Vڥ���[xBgѝE�a��u�)4�H8qm� �\�$�y���)�!����a�)x�?��wEcȢ�o�~m�baPGv��� �⍣d��9�����x.^b�G���j�6I��s�^�0r7��}M�.Bv +� ���m54��dL�ǶVJ��8����^]_v9M�i�=G���[���H���:f�s���>�<yV	�=�=q�T�t�D�ʕB�o�`@v��,�͝��>s�#�-�Z�N����`�Bx4;P>�'/-��"gs�W`w���+�w����g��E��e@]�O����rb���0�s`�x�T���Ch=3�Q�����S��`e1G��уQk��k{����-I�t���Ԋ	��T�|����Q������d֐A^
��)aЋ�$v�ٱ�ٙ�W������bY	��b�f����O�� �`�8lC�pa���w��rq�8�{w��e�zV��F�ͽ���Uj��p`l-��?�Ũ�(�Uvq?H*����N����b�����2c u��Mt��{�s���.��7l���\�� �\_C��w���
�P����K =��XR|�}��c������K�����|��H�x�pH~b�%��<�����s�/���8�|GiǓ<�����ϭbiǅ���#-�?�)Bl��Ip6��V'p��]A����=5�S�䫱ے�-��muoʣ��Ư{*jڢ�:������w֌<$�� �9<F1���i� �C�"��lR�6z��^�o���-K���`3˼V���3بy9��ɥ�p�����2\�OOl=�:9��l͸��ͱ�%�)GsWc�S�ӽ������p9���(����a6^�`�=G.����*?/�����:��B�:�����H�H��1������Jr�u���I���U:U2wx�!������.9�1%G�^�(�(n/�
�n���8�- y�kQ�LO����l3y��{T
����KF�5�'UO�A�ԔN�A顓y��&2�Q�-��ŊdP�[魙_���w갠4����ץ��s�^pVr�n�S>y?�T,�i�� #;��H%�R��rT��,�k���?�}�і};!9#�]�u�^ ����u�!7gA%�T�\���͕{���B|v&���mI��ao�گ�qm�_��9(��K�_]%�$��w�޸��F����V���cL�P��kM(�n]�1Y��{ظ($���<�,_-KI���b�cC?V>���Z�*����nfCը]R�Z����՗�Nin�����BEi��'½i����D�.�d%I��<�3z�d|���إ,����EqP�b��6�Еmp/�E�Q��+#��k=��3�.� ��U�������N�V�{�+ҥ�WV����z��0ô��m�<;��Җ�t��s��ʿht��b���b���g�8Sj��޲��{,���o�$�I[�zL����n����C�%o>R}���g�,��]tXvtZ�����W��7�Rs���FKw`'V�u��3�z��慼R�\�K4L�󬧇0��`gHA�}�9�ٻr�7��+�E�)�1�rޥ��B�&�[�G��C`*�=&��2�M�C�L��	i..iaߘ�P��'��y��J*���;f�ޞ��Mmp�����	�P�-ɠ�g��!�� ��3:�������+#���������x�x�ݟ�Í'ȡ�̼��}�T��9[O�����-b�&܏�G��V�����@*&t��J�_��[j��qG��&������(f��5�s<w|-�R���f.�?�A�pvl̠ p �g�P"�3_I+9��d~Q@�u-�ʧ/B�pZ8�5{QN�SN�v���bE�8�I9O���I]�;u�ݎ|� ~���Ous]�A�=�h��5������*��cN�-Z(������t�J�}/�ֺ���2,�M����4J ���8��53���3`�A���c0�恻��`�ZP��C�I{i"������8V��v� �~�^�-������C��N����@�Mo���w�v����iϬ(n������&�Q�Q2�@�X����D�,
��q9"�M`�6�M�@�f�߈��K�+Z�џ�T`�+���y���a'��FK�5]�7x��n*�6���t�3s�뒶E(�Z.9����]Q�0W�����\��÷����0��u�BBc��_��4h?�⑓g�u���<�+`>�:�늸.?bk^�~�y�Oz/�G� I|$*�^��H`��Fm)��7˻�P�#:�7�9vM��S��FO@���~e�$���Ij�*w���Po���~o�V��|���0f�F�S�����,���8g�ơGy��#���j�~a3�N
Ā=ے��*��ǋ~]��:`�M���@i
ak��d��$��h������9�_���4���|��,T�U���#�)D/Cه�|�V78���qn�Q���+.:��V�hd2���f�W��@ K���>������n�g��qwu:��$�.���	�<@��4�⌱��b�JǇH��-+_��GN��.ˢށ���z�"V߰v&oB����8�낌��s�BqȀ)����ª�H#78pal�K�k24��]�IK0�.��=�*�PxQ��{ۿ}�h�wE��d|?����*�s��zA6�;�@�ފ'�x��M�o��t�;�^'J�k(�!Lĕ��Z�`���%�2ׯ��y_�I�^y�����z���4C��ۈ�����&���>\�+`��}Y�܃�������ӸT^�X�P�'�j�$�����)�dJfK4�Lbo{�� �M�櫧u�(�ӂ��`av"4ou� �VF�8��=�V�Dx��x^���B]D���7*m6�|�{;٫N�C�?������CE�5��"���#|A"�(U�=\��ޘ�V�a+[\���K�F�x�;���6�~UHy����]4ͭ�?��ǢtgԶQ��O)nt���W�U3�=��M��(���]Y��TO`�lt{_��O:Z�b[2`FCe�=L"5^�����sV:7�,=�YfLNe%^M2���Q�o/�n� �F�.*U�F�ڀ-l�o��A���<�$Ճ߹���^�6NLk \}��Z+��.�m��r��D���d����I+�8�� �n����Z
nO)��z-�+���Y���[�[JB\�l��p�R�G��
Eu�)\
�V�y"��3i����9��
�7������U�EC�/�(�<��ʩl�PtQ%�N@��t4IH,*�
�79����~�3_D8/3�".���4��`�e��S� �����ZQl
��j�ө��o�R�b�S%|$|�ñSx.&��I�(~ �����\��y�-j���k.~{}��/���E,�C�(N�kt�������w��Q#YRwp3I�N8�x:�,�i,M�	D��T�Qk�ç��)M�D�(�]Y2~,�b�3��tS#��9�00�xD�%p��ｚ�o.0��Q/�r��a3
v��g��&KXb������ȣ��l��| rO>�.mY���f���jfɒ��¿>D �ֹ�S���G���CWմ�D���
%,e���=������B��s�ֺ�XbYԢ��yT'��Xă3C�Gv���hYT��4�#�yu�~��{�h��bN�O��p�;;�8�~��[?>�q�\�<AV���4�D���KMm8͂>�3��y+�x�җ���^T��}��p�9�b�7�-�C{:���46Ж�7&C>5mg�������1�)�U�WLQv�HF����.)�$��U-��Tqq��ި�Ǡ ��!�b߲�S��z���`��TMI�8od
j+;�2|���
9��<P�b�A��Z`��Y�@�o�w�2�=�k�q���8��Uk�� cR/{U g�� �{'L�ec�*�	���k�	��n��w��{���05D}��X�~��kنzVE��7�HM"��P<�"7��,()݄�VTl�a��u�����U�N>��"{}Y"������꺹�%��4�Z�d~��:1#�'�OJ���}���1���h"�l��m�����w&���]Xr�H��n2�8���wO�iOn��-A�Ǔ�r�Z�@�V�R��^'7�W�m��kW|�J>mT�C� ������tЛ}��㍽&*{��HD�dcQ��s�J��gY�'���NȚ
��Ǟ%��co@C���
DT���͈��s�����@	3&ʩߨ�a�R��j�<~�(��\*	\�Qo��λ�61�5�+V(�r*�U^Lyw��"C��|�Eb�+����o���|4�@���H �'H�Η?\��U<��3Ụ�+��T�@=�[�����G�u�y羛i�	��y'G@9�g�X��c�ߗВ��]Ȝ_%��М8\�����KS�G!i:N?.PF#y���͢
��T��D>:���BUcͅ�o:��@�\�x	ԯ�����fD��L����W1p�ntY"`���#���T�jP�h�O�8Z�U�JX��oczg�U[���6x>�=�bu���d��' |��)�)�fA����Å�z�v�jWd }w:���|y���|(�*R(��mm�[18�� ;�LXS�#y�Q�'J
���3��2�1��Յ��J�+y��B{����}��
A��o�⃾��8M��va�K��}��J=�@�6F�U�Z�=y�3j�*;��)�N{R�7���0�x]#�dS^i�y�{#�8pn���P4��R6u4���ǻK�f��!����#s.���ͥ��aG�(�`�u��j��g8��y�Kq.n�����A�c��������lcux@�k��">�����7�tмy(s;d��4�ŴbM��N��s4���E,_���i��_Z�������*ĤJ�U\��w!���y�6R�|�|�9Fؐv�A�b�[�n�A�WiT������_�TO�e�#a��_.But�[����t��g��~��k�zgM���D�Jq$%9i���$h�ul*���j����v���]�\��o_�w��*�#��O��4rfF.v�j���B)ʑu�8��=*u�����Y^��M0�rapK���X|wA���޶��Xӝ��Ԛ`LSS9bP��]20G�CϦ�b�Ju=��q��<Y;������j���y���5�L�~�o��л�|���\��&>B��Gy�<�ˣ/$l�v����K1vg��j���7�n煌DIKʲ�<�Z���6񢎣\�y9�"�K��}ZU���\C���V������������"`oZ��Q�qoC�.��*[-��ef�ȱb�u3tR���ue�Au�iU��&fe���A�ʤ%X�	���s�4wT�A��R��6p�-���C�3���I|����~��iϋ+�V喀�+���w%����Jib/X�Us�óU�(|t\�G�ӽg`�!�8^��8_�z�x�փ����W[��'��:�.���.b�c�f�(��*��ږ�^-����L��Sʆdg�~Vy��p�C���tDf�o� 	q$�	�iypZ:\v]���ޟ��0��7��^�5��YO�%�����wxa�Ǽ�ag�Br�n�Dl��NI�y]�� �EX�d�j�l
�yH��I�S\_��ݻ;������$�����)��^�9�,' GCP�T,��ҭRo�|�ڱ ����򷹕<o��!+9�P#�����fǴ#���qty�.� ;�뚧�
��e�����<��k���l��F�[�������M�v�A)��(��طTv,7J�0vXh�t�y�.+�3����2�:��p��ڐ�|m��Gzp�d�q�:�����9����1P�D�5a�:�a���w�|��s߅�����Z�r�ǌ:`�&}Qp3O�z�|^�25� �1�C�^�& (6�x�v:ߴp��ƚր������	c*�_��G&;e<\�j"�V߽��w�~�죚we��G9�n�e�-�A�{�U���(����X]Y��]+^�I>��9�7��=��`R*���V�#ٓ�~N����*)�bnpb�>��ݴt ����[�H�|w��wG���F�5��oa��t��4�li������og� e�*o���H��A0k+�o�]�޾�q������^a{L-W��c@�@7O+��������:�t��?Ot�U�B�v�G�+ �9��J�����nw�grת��_�;x�P��z�1
��]���h=��[w����)D�A�p(���wC0ds���9��>�k�F��Ȫ����A$�k	ox_O0gT2��3��6�~ƨf�s����MN�s����ަ�t+���)+�yk�Pʂ2օZ:��^�S]=����:Bl/(�hq��k'�{6���0?�p��V�x<�@����i�}��!�L��G韉��g��l��i%���B�:�r�q��