-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uwpypXiF39l9xgFKmqReNX7c59NZbf6hf6R51Us0eCuAMSBjECDBV6chBDSVxoR+Qvz9mCBJ5t+c
lT5/3W1kLavvkUVnXgfATL0wOCOqtZdILY9O6if6I5AzHUFLvV8e5zGg1Fs9IK+OderqPN4UxzU6
xaWgSOdQRNRpNrfoXymrbuk25Rw8pzXKOGwt6B9FbSDz83xgFOMd+e0f+D9qxPXge/c7tvJNxMQv
qCuZudLjfD87gwQKHTgZHNJDKolkygt2tXm8jv7J/Cj1FvRkwJ1sKYpuqlZ3vjHxPp8vO2WRhH3C
SbN6Tr00QTq9oaH5096ayGfIYwyL+yOnX1Phjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
nhbHQGbHV+HaQ5bPD4js1NY3KLuxhkHS5ToUH4Et+5JJaCW1IoC+G7y48SBci0qZiv6hcr2bp1Fs
D1d4R2ae4DQFtZuFsiRYYazjnMv8iAaJqKJO2A0UfhkAfu6Foav0aK1+9KrIT94NgmisIO+eoh1K
2VtSkZEXGrs1l1h7SRDI0uVS1f/Q+fa6O8SSQ8Lm61FMe3VUn97gbL1rncuRKPPyx+dlfIuVGJpn
JcQlOW3krx9kQgtI/pXpN/0yYreIwWNa5JmKphWUMVPay7weA0SNp1eCR1cqa+fzsKtliAi2oXXA
llLmtpM16SxVY5gtvuS7BHhxlXM84dTo1xkcy9nWlbv0Zq+VqzdyTAVKOOwTy076EPtb7v5r4DH/
a31HTTA1kthUd98hMkwaLoK1+uFPEI0myejfxhPv1wL25jUNEhT2FkS8+9AAcPk/WcJE2fI53zaq
PdGalThQUmOIUZDUbIYWiG+qII4zuAtmLYMAaIuG2pcNZQoLec1bp/nr7rjWJ/AAKT/gZAnxEpe3
VQX3Ef5+QpLz4t/R3xDYnF8KA1xQQgpeQejXUPWGmeAvcRw/2QZy3REZba4ntSzRh/dy2NQDBe1n
vi2Rz+h+/65MeGm6eSRkDNdeV1dkexT+8OMgmmbeG+EZ5IiaE9f4QTr2+49ZRUfGWZTxjIEN1Xnh
iNu8deui3fJa/q7GX3XHkv9xuwlaW7uaOWFolJM6iAenBikzaqwDynzPCrY3HQz+36Z8tSs2bf56
vSts4LzF0qoq0O+Cemd4VQR1RtJqIlksoxHxuQR2H1ncxJ7NhUDL7EDsRe1LbCC8LANBUid1dSU6
/ANpWkk5lCIkD2YKoy9ZouGrv+KbfuXuwjBr4C7oGn5WMIhnP6//M2IBlUcF89sS7fbbOnImbiGU
V8TCMUXrkE5/D01qE0jx/cEWfZWjaeArkS/MpB7Tk0ADX1TUjXQcSzrxPWpJJxHml776HuTlG3Le
P3sEtP2Bd42qzOL+xOndzHLqt99s/52Zc/Gcr8zppL73fAi6/Csecy7TmPYVZXkiwzUbfQfvtrz1
nrzXb94EoxwVlaTS1urUtYNhfMqbcd2SaqpE2hhQTpjtButQa550RuMuZtOVaDTs+/F+h1DIlDKS
GFymmeXwUlxgZLpiUJZiWEzTBKTPH8XGpe4WBoelWsXJA1tUwHGsU8XRP9Q3RvqKrtvBS8kYf1LH
VFnKdsUgD76RCulYuFY8/2jAurFiXF9Dli5rSMZusoEDw/K/r9kCV7DuIO0Naemv5BEQ+hmAvADj
Jgp1Uc+0pS9rMlktEfYwsfwZL6w2C3hgb+8jGnaBgMG7k5cOMjsIMqJgi5FPEScueNdBw4y8DXMV
1PqUVzzZx8jiT13RTZeORKqLokBhobRDTY6lsm6d
`protect end_protected
