��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U}�Rtq�O/h)�# ��	��|�bi���$+���>$s0�jtڭ'�M� �b3gC[��{�]Z.&#�s�l��@�Uw4�|DZZ�9S,P�È�bF%q�k`�.6�BX�y�O�?P#1��h=��ҳ��������Gܯx�!��=�R
(7F� �I�Uldc-%��+t�!��5�Y3�#e�$�At��Ѓ�nN�{�_䟌{5�b�q�@N��*�{�����c�-�w� 9_Ԡ[�H����/���	�O�=l��e�<3%��>�tɞw�Rҍ��z��ME~)���mpo˱KX��[�sq�q� ӥ�u)�?�@W��K6DcW���zU�=���륦�� ���b0��$UL���gq����Vu��F�}�l���Gk����WY��)��A(���K�L#Gg?� if��l+�_�&��No�6�G��M΃�In���[�[pE�����c�m�k�,�H���
��v�WVO�2���J����`�MLip��U䅣`���s3s���#t�e�m_�'ܞ�"K��2|P��-��r�c`��1O��P���}1	E:�.T�v,ʁ˯vFl(�4dh����jtc,�����>6�VX]�>V��IM =��Fhs!���"鰑����e���ѬBEU��U2;�'��b��c�~��TB�*�u ;��(���k��/
�X�eV�h��vI�EN
��܇z��W����1���ء��{/%oZ�R(����'o!�Ƀ�xT��}s8��&ֿQhU���=�"�L�醆���W�?��:z8/��0�f>�����V\e�ԓ�۪���@�����Z�\o7��ae%�N:�ځ{��O��.
`���	e;��{�v�����ͣ�g��e'w���{�z�ɦx�`�J��+�Wϕt�X2��b��ʛb�z*�����+�&��_ɤ{�h+�^!~�so��!C~������	��f�I��P%��AA�4�'(�r�'�*���5�ٰ]�:�������#�ѝwx"�I�Hpʞ�8�GoaLA �����U�x�A��<��[3��˦+�؊q����/�C�Ģ���,=�~?��!x�2i�I"L��3���tՏ[W�O���c{�W���N�S�V8��!��qq��C�E�Iv�Ax.؋�<�)�X�Q֒y�݃8R��?�k�liq�o�����>}A�TܣIODv��e%߹9�.�0�|��04��aC��kj<��S��{5�Z����-�鍷�CH�j���T4�S����	�(��NV��(F-��T�آ˛N^7>�Ἦ�G�X��ļ�Қ���E󙷢q��_�'�rqE��^.�X@�:�����̰�O;�z�(�(ܙ��u�f�Ig���ѡ��a[�ka��J=����'!��[4{�ڔ4"0��L2"9��\2|�Q����aOnjn�,f���Y���p���.�D|D�ӄ;�*�)s��5+Ժ�Ȱ'����?x������/�ݶu��!m�v�@��[+�p}��)1�A���k����dgZ��0pB���'���c�"�TÁ�<�S���R>��4�>m��K�8>��Pf��^��%�	�j(�p��#�dD8'J��i�X��7��
�S˹�$�-n�*��a�.��E[�����d��� l���-�5ɂ!���d3�ə��><4���p���m�T��Ao��cH*M^�����4G���y����}	�k��3RU�:�p`���,i���LP�{*���
��Nq�u!�m~��tbr���k�&=�o	��Oe(5�h��ȧ�W5������Fu�#"GĜ����}xp��H�fAN�RI���@D�Ǫ�.P�,_�8G)�-08�>�uGF�������Cj�D�Dc�w
`�U��A?x�L��5$Fm1��3Y9��i�L���M����Y�C���+�d�zsV_/)���[��;u���/5�nK��5���_�\��L˸�=܊��m�'��p|\���5����r�霩�Ǫi�(hf�!'@%���L��B3��^y}*$G4t�Ot��T�\=�2w�z#%�麘���;�e�9׆�\�.�S�����lw��a�jj*&9�����������,�*���|�_%��K38M�wC$�k��K
�t2�^��6)��ѠAz���`��Kk�4M��J�^����ZDZ:�S���}�SG�E���ةP��/8�;�7��t67�߿�(h!�귋��g��UNù��gv�%��d)������ȩ����Nɐ������C�1�����06KC{+
�����4��I��}j
T�a������T �Oo�i�
P{������@��` ��T���u���n�����+Zѵf��`Ǔ����gͻ���?Ԋ�Mc�v)/�.}��ݟ�+�"s�y��5������yT>y+3���i�H�A�/��~���TE�&��6s�y��P�i��!�2d�ရ��S�z:�z�.����#���r�dܛV�D2��y?׳#a�xt4!��A�#�t%�����|s-�Q��]52�4q���X��y��â;䢽���wY�C��{x�X2(���`mT��?��; �(�
/n����D���K��j0/����
W�����l�"���lX�x���q
���k��S���_-�꽽k4� ������y�祒j���8'̯���6����`�)��Q���4�>��?@��>�RV�?=�H0	ϮoS?��%�&Q�:�HQ]e�� M����a-����s:���qҼ�
���ܴ�'#���i�b�	/掚���W���?8��!p�*�w�K�xs(q 5���sU�H���{�����A�0i(�g��-X�W|�1��k�)�܎��T����Y�\�M���Gh����2[�<���K�Է&�q�W��)!��罭=eť>y���F�o�R���ؑW�C�S~>����?�z���X��k����̱7f.�jg�g�LF�5��?�Nwz�����b��i��I6�:����l�Iu��A�o{zP�m+r��i=������`BQTҕj����a��:\gZ:���ӓ�T �������E�J�wLWv��q���~�"ny�ʊ�ԭ����MܚqK�dX�\_�{�z����"���{�'ێ�v���1�l��h9��`�F����hU��b�s�,���;��)�r�k�Ə�/�%����j�W.:?��&5`;K�,J;8O[�{�����P�0�@���IbmS�ϡ�V� �+|��\�	��L�9 �_��O�v�:0��m�-*��.�3Q�]�|��_/ts �vQ�>/w�B��D�XTc�z=�3��3��:wL�ɔ��/�7��ӃVj`u!�x��+'�n�,����K��_�
����������q�%��]-�BG�Œ苋O�B���D����=����DfS�gV:wq���U�F�!7!�,UI!�0i�M�d�$�Br���� �\.P�t������+��d�4�u�VY���	�r�D�n�%<�7 9�G�y��I/J&�:�ӝ��]e��z��r����H���er�+5�}�ż��x��V������N��" ]�'���|�$���;;B�X�f2M����f��a"A�D\��}�%�E�ʉ}�� ��O͚l�E��	�D���IX~�YlO��L��1i��\<Hj�
U��ϾQ���u>�*��� S���K�[=`�JjC����N �j�/�G[}D�X�	
��R��m�	|��ru3ZY#)��~�#ɫ�e�r&2i��8!2IeJ��0�1�D��ԞJ���JT�?3�xWW����;����d��{��x�mQd�����Y��:��Ce_�9�ХX�ڼ�q���R~m=&<,E2-�3l~��,��p`���Q-6�Ӧ�F���5Tbz���}qgӑQ�1���KP4R&f#3}e[H�Y:�J�@���4���r���7a+N�O�ò�P�R�I.|�G�V&"�����~dB�JS�$������y��B]�/�o;���D��x�{W�	ǝ%�>_X.�l�?�
��KE'�R�&��n��H��.���/�r��a���z�� (�� Y?�1iw*D=��Us2�P�	,��%>A��o��9���G��[��[8s牛a?%���S,���<�&���%:`��jq6�ᖭ?ZG�V*���3�*�$�K���?��.��\Ģt_��H�b*�6����o�;�����V^zͦ�k�RWcI]	0��_6�ci�gYu��7(�y�l��6�߬d�$uRj��0���6zA�ic��dF������r�~z;�ӱ�}�����É;t�/�"���pPnJ���ԋ��Il@ý�_\��~��tA�qx�C�yQ�7�{΃ٹ��
h�宷maH�ݕ��Wqٱؤ��J&p1�����%7�?y�P|�o���
�#	g Վ~7/��]�k+%8�c���zn%C�.�'!C��F29[k%�e�*���zCK����;�h��,A��S7y����~�@
��󀤯��Vf)J4��nj5��Q;`v����=�r���!��m瓬�5��qp�)]�3�#�$&����G(I�( ��=��'� �����i�,bg���L���w�#�7��핮�V;s����V�U�J^�iRbx͌0�O<%Y+o���`�}b��5b۽���؍�l�6{��$W{3�|�<<¤_�RZb �|�v�"��	��5m�3y����o5�@��.H�.����(⾁����*�f���=?�+,��n����1DΨ�:.8֎�\������O��:������/�i����L�2K�P��rzI�줣,��y��S�t~1#��0����<~h:���;��/4�mI:Nz�dy��n���Q"]ʰP�r����[�m3��6q��T��p0�
�O��k�)#`i�ⱻ�!I�<��[.f����Ôf�X�&�����\�#��?�c����uI�.�N��U4�O� V�h�k �E�(�"R	�m�^�Z�@h#}A�H���)/��*&�~!�(�ՠZ��M_C�8��ZWx�j�ƶ0���fAI\d�ݽs���
��f ��/Mf�"h�g&ʿ�i$��H���KĬ#(M�[b������W�&��,�`�*t\���R�U�z����X ���5�#�E٥de�kR�T��\�x+_� h����!�"N҅U�/K�j>��'Vin#�M]���A�C����럘��(]v5D}��l~��伉Z��H��ul��u���~��}除(�k��_0W�A]��nc[�	�J�XY��+�w�xi�a�P��h��㻠��?�" փ�ET���;.�����1�7�F�#/,�#z�>K�ޏ�X,y�t�����ٱS#gx����xKW�)Ҩ��e��2�6�M����7�������fX�Rz�p)���&�ݴ^ښ���Y��T��*<���]�75Pq���ZʍqY�_��QD��E<M��v�0��#����������n��񦅝4)�G�����s[kpJ�=B/c$sG���-ET߆>U�~� &��3[���z����-^�믇�,�eq����q�R.�d�b����:�+�,�3���qC�-9"O�G��K��ؗ�+��'�+V���?/n�a���r[�{�<T�:Vdz1Ɏ��J��ɤcl����(�U;�R����˅+��9�6�]����ɒm��H%��f\��(yża�|�W�i�=��'��|�t�� :�����" ��X�Q�"h����	,�k��N���)���#q���`I�)�,6��O~Ѳ���<u�h�\���Wɗ�?@���c{4oj�ڂ�c v((��͡�ՠ��_�!�_������s��7�CZ�0T;�/,>��j�t6!o��dMd��!<X�֋��:�/Ʀm�b(�e��b��e�(P�+���Ȕ�@tl�c0 �yK!^-��z�ɭ��=K�t����p�0�ָ;�%���:MU���\J_C|�!ݲ�ޑ~&���	 7�KTI8�z��9#�Bd��OU�`;���7He�2� *o�f�|��I��d�"CHf�켱V*��������B!B��Y�&U�Co!���S���z�>���5#�Z�ɉkQ���Pܩx)Me,�ܞ�*i��C��W�<�o]�-����XIu��; +�.�ٟ��(��u!ܞ�E��bD�[���RWh�mçr�����>��h�
��D�F�6�+�+Fb*������b]�)O�S5M�jT�5�'�m;�A�����'I���|�x�DK̙z����ú��6�*�i���9S��%m�6����B�c������]��&&���i���/�ab��Ŕ"�'D����k� �ϐ�k� w�һ��<��{;��&��}ޫ���p;FN
�s���2C&��y�ꑐ���� ���.<>cMZ_2���H���p*؋E!�U��t;'��$�TU�kό�<��oi�i��n�|�c�T�1������J;6����1�d%2'�\f���z�*Y2�\�!V�++{��|�1�B�F
�R�8�����z��Ay��䆐���"o�k��b�z�#�&����7����~�]ƗfjI��o0�f8 Y����fעj��AJ<���Q��;Ұռ&wm��S���L|eLX��l��4�&���?�;���낡.��h�W��?i�F}��K%R�W��s\��[�0�w/��0@��WȮ���fdMD%�����Z�:�~�X��0����H`�h�h�}�*~a��Xt�V��0��r��m�;T:��x����fN����t�@�v��U��Rb8_χNw����B������v���\=[J� M
ټ ]%��y�.���g�)�VG��dS��E���\��[b�N��۶s�r����I~Z�0<`^JT���6-��k�Y��L�V��}��R߿�=���!�T(!�%9&��{Q���rP��?1�%��Q�<u�R`����g(r���mWt'�/<yK�#l�X�Y6��h���'�v%yQ j~x�li +DxT��C�n��I^O*H�����'���W�|̴�<9cw�IF�Y�J̏`_O�U�L���8��؜�~#�u��0@\�xe�7�u� 1�J�dp���BBl�su��9�H�/O�p�Ea.�nW�\�3kd�UDR�O���k�3k����KX�����U'}`ה��$��B6�Ed��(!5�hl��/)��_܂�=�*%A�%p�0K$��V����Y2%�Y'K|7;�EP�~��L�ٶ��t�ubŴ����Qbc����`���8'�F~�#ޯ%��^�6ԍC�ʳ%��$%�[,�ePz���
E	Vh�+!��'2�H���X8��?��yQkq2V���9�qQ3�R�$}�X���l�C��F�)9&�/Y`��fȝ���f����6�U��Åu�ȟͪ��]H��O�<&��I~�e��ws����w���� 㙫�J���
��X�M^{d��칏�}[]��I��ݭ\�A��T�Vm�*P�I|vafok��\�nI�L���%X�l�&�y�(�,)8Zt��
I!���W{�Z�}6�����Vt9ܳG�7UG�`ې�ک�#�;�s ��H��+B��@�AT�Zf�(���s�#����s�z�"Ȕ�"07"��ٶ7�����̳���4��	Y������]��HX�x�:�K��j`�M&^�X�������$p���?/(��'"�[��ڳ�AZ ~��(Tg��~�oG���!�㼤l`�
�N���)�'��ǯ��*�?BO������ՕF���֢��K��F~���Mmwt}�0�+M��(�z?��@�4�b�
88�+����r����o�7]ʕ�cAc�Tx�]�lN�͚O�]b �w�� |">/rQʥ�Y%�2���b��$q�l=��T#���pfݥ�f ��� hF��ܭ����7n��Q�U��X�@J�b~�s�Zn�t����4<)L�Gq��0�D֭����v<c�[%��S>A�D ̍����PB.�u@H`�z5�����nbbx�0Sm�p`T(�w!�
7@~�'j&��� �ɹ��J��AS:p"�]����=@*q�	4����n�����CL���M�W�v�{0tc�����{� �!��+=��ۦ���L�)_���$������F�]���[iYX��U~��\H�����Aёx�Mn��uuM>�b�*P�eH�Qu�R����a���:��ٝ�-hJ�(�=016��דŏ�7�b�X����BjK&��c1&q�I�A��E��=F�N�����gk����Sl�	�-uЦ�
ېVǉV�0��[.�NO��;̷�L�`������}~�:�>��f�P�"h%�:S�v�C}�c|��V�<�D����(?�9�Lgϝ[v�݇�P�N+~W���Mܸ�������1��A�������|�/�g���\o�������/@�q�hnB��@�dB5��7!�"�+ܷ�zl��B���W��r��a�A�o��x+i��!'[�@s4͗M�j	�����۲V$�s�����k�YB��K3����/���k�m��oW����)�V�[��i杙����X�����飾&��4�~\9w����Z�	���M➪�t� Z��}T�ܡ��x���Ί���/�h,Qp�<��3}gj���O�-0�2)�:Ƿ�w�9�{b؃.e���|H�R�(W)��v��C�h5��U<F��p�<R����(�yo���1^J��<.In�>�e̽�^)�.!=���@C1��D���������H�RU���"m�KQ�Ɇ�wA�S]?�cN���L/o$�-��z�h���t[l�a��m\$����<���8�Ӥ#.�	�\6�7q�������E��@����#�ij-�+�e�6���fJj��P/�vV��_�" �y=���0��-�[���\�k
�#��S�=�/�w�j��ϊ᣾^n�-'�ϊW�`�y{@��B��ܥ��F?��~���6%��5�rq�z�6
�]<l��kr�����`$�5:M_��+r�?�zw�����8'cPF��U�h��p��"Q���rC~� 2��G�F�.e=�����ϋڰ�|�z]L�s���0~��#�f�ʾ��b������[�l���x{����ڄ_?8Ȫ\��!�0�`�7p&@e-Eӈ����v�>�>z�$dz��fO�g}����`�<NWކ��KYƌ���4����E��z��X�[�����g��|K���^B���b���e�s�g��~q'�M OZn�=���t��Lt�s �S`UT�y�Z�'����D�N���q���&���_�j-:^�ֳt���81���������4���(u�L���g��ɭ�mhb���k&�Q�Jc��ن�m�Q9�\��گ��c ����������*�l퐘M�sj�׃�{{�P� ��}�V�YI�T�@��Ƀ�!�ޣjaP�R��Y���r�G��	��byo�a��'3�3���a��|�=s�\���w�D�l�+a�Z2x��r�������:����t�u�a���.����
�����XQ%F6�k?�ո�͵c[Վ��W��8���cs���DXn���[۫�� 4?��xxΚ������5�v��6m���9�`����C�᝹ݕA��7��y��$�KN�g�ގ�O�` �PУ�0��C�����[	E�ڛj�Lݸ�9ϗ��qc�c0�[�d��$v����'B8��0/��Xx���=OWa]���Z	�M��o���lqZQ�tCNVF���扇1
����CԼ�Է���X-,��ȓAn�8
)�,�?,�����@�/�����lB�<NȢ�����r2��o�q�E��Yb�����I�$��Nm��!�T���`��T#1�J���b�d��<��a� ���ϴ��� }c�gk��=�/��@�8���$���.�})�K�]�X�6�3�r'�p���O���#YI�~�K4�^�O��h;��|s�?�j�>ň��� /�\F�v�E+����ID�d���A���Ze���]��v.Dr�%EL:&J=7%`���M~v����F���ތ�G������~��ޙ)�}��X����2$�c� K�FO�K;��e�ʞA���2��cM]��4�ݷ$x!��1�K�P^�I�7�?	ʿ��ւS��@�^�sW642N""���'<����doGHB�������ZKQ��'6�M�L3�&�Ɨ�u�b(}=��F���O��i�9r>F뇺[g{�_�<ә����F�c�	�a��� Mf� -��;"Ņ�"~���ዿz�a���ov�~����T�m�^A�?9{֕����F�I ���e�i��CIǀ���gsD�'���^©�3��֙��Έsj4��V�-k���_X�r^(q�~?�).�� *�nm���~-g �8��p���=�=!I?��QK��^�nw#�H{{�y!�����E����_������}�`5�1����揨��w��\���3�1�.�;�˱��s�m^���"Yt�2��D�k��Q7�}~ǅ�Pݯ U5���{0'<r�4�\{�c0�Gw�Q-\ygo��3��_�gNOZ�C>���#MqnN�dpn��Y��$�5�����+��(��`�u�>��,�cl/n��$d	�os3�ł����λ"��@��c�9[ۉ��H��ǡ�W�9���l6����ʬ�}h,7��8J���cD{�L=�D���_�bS	6�/Px�����a�D���c�[���Xi@^w�i�	���s^L�5J���e:~lT<�ZS�I�<�v{G�����9�F;Nv΍
��Y���㑅�`%��ԻxA{����N\�=_��|��	������"m��~0�Ӽ��p"}+��[�p���bb�)1tʰd�~�Z�\���ݹ��s����W�l�_рV�@�������pd�X����)�e���=8�A�2R���q�u� m�m��wȅlSsQԪ�D�겿�.���+�g��S�ĕC��v_a<�´Q *�����n�I��O��&���F+���b��-��$���s8o6�t��h�+�� !�f�A���)�7A��T�d�D��\�UYy(:!���۶����ᆪfꃐ��8�v�
�\8;`��s8�5�
D~�7CXXْ`�N
�>=��wN���4�܋�ѿd}/�=#|ER*��\.,�V�)���$S(�Sx���G�0�ߖv;�Z�I�"*U}��1[;J7��Dd�B>b�h& `#g�����r�f��BP	���_��+-(> 
���n�����uT,#y��jA$,�>{ɣ�U�"���� @#��myl�(�����y�����r�����8|���s��D��o*o'[0����[v�K%�X����J��Ǽ�@��^s�9s�\Uvϼ/�[K�6b���T/|-�����\ꋱƶ�W�ET�m����q0n�����rWG��Ō�ɾ��>�����n>���"H9�w��ڟ¾���@o,-LZNs��D��c���]~�nH���߬���G���6��Y�:���%���Q��R��h��x�[|��%9���H��^i��
� �2�;{��[�M���~���}gI�M��9a���{y�1'X eN�0��˜� ��D6�6��
Ɖ�m�+�$.3���"[���rlKc4��
�{���߈�Gx'�6��ô}���=�u,��?�>}\Iq�=^I��6��*LɗL[l/��k�}�b�SG�5ђ��%+}eg���Ic|�;��c�6X�׮%OoHR��/�IJ�Q4�F���y�߻cs53��93�x��z=/f�����4��$��������O�O
nޭ!���-���L�X-1�}�kuL�D�`�m2jR����:9��z�y5�սrN���)6l����{e�m
�7�r�[�>��Pk;��]����"�3��vD��-��{̹S$�XՕ׹�:�Nf���q2_��Lov���/2����A�TY����b�8�	�ڞ�j�-�)���IՕZ� ���Ai�Kʏ�
��j���*�ԅi�?�S:�6���L3/{?L­�<�Qn�"'���A�l�O���t�i��7d�At�]��hID���g<fҵD�?�Pm��Hyq���n��*��:&wL�S7s�Vc�2پu�T��"�+�H���uE1n�u	���(-�W�-��MJ�'4Ѕ�a�q9?i\@��8�NL��0,�p�!;�Q���~f~�I�nh�˛?7e�VK6yص��g)fY�����&mF���J\F�>�_z8-�-y6&6�&F�z�	eB�Ӗ|�U,6��~��䅇(�+r�M��j��������;	���`E�2�6�`Wڭ��q��e���ϒ��t[9�4gN��f���0�"σ{nVRS�Yc聬��ez�C��tp�f�(�W=0�3DU�H����ؒÄ"�Ĵ`���AR��r.������S�n��G�Ox�>�\�/s���W��k����o�ᐲ��c���5i8�cF��z�0�v���3��sCC��w�� �,i�s6G�ecc��̈́��$��V���B�d�YFK� ���52L��a[փ�\����
z͈��c}��{G�,�e�b�[�-�7}l�gi=�&��f��}'�/2e�n��4����'������%�� ����0u|���������$�2oΥ=v�=~�2r���ݒ2K�;*P�Z���2��D��P`H�t��{C��]LprD#��Ψħ=S21��!�C�o>�f!����_�)����Z���Aͅ@�ZФ3��&�1�cT�&�Z��վҒ�?�DFq��e�̤���S�ɑ�3/7}؈Q��*�"BI�y�Qo��,a�7�k�b��^0pC�{!d��3@]�� ���W!b�a,GI�a�Iu'�w��?-a睅�T�X��3�2䙢���Q.:79�<{lb��M^�v!��u��ϝ��QY��;=dj^�H�j�H���b�;`;���eH�8���4���ճ�x��l:k���h���ZW��<S3���Z��!�F�AV,��)~���75��Q�͢�G��7ڛ|U��/]F�mQ��'_���.U�zo%�Αl�i_�_��Ӥ��a�_K��B�������i.g�s����㩍�J��b� �s~Ջ�� ��*E�v�"�@G�0�؁�_zi��	\�8�(��Ǡ��7P��K��<?�xi�bW�7��t.;�q1��jq�
� L?�7����Yx�(��@#�>�H�,�Z�k����dQ��矣�/�o�:/�癝槎��v��f/�U����F��m��ϰ�*��B:���;���A��[����9|�9B	ۂ0���o�҄�:����@Q�8pWHn�27�����X��P=c`i��\���R*���}"x?�B�V��Hg��+D�
�y���=��܀\$�n�ٰ�PU�S� �t`�}��o.���48Z.0e��Vڝu���җ?��$���-�K o5[l\�UC ���`$�.����1e���P)�L:���D���hàA��i}�t���\�\�����WB5a��_��+E�
3��R�� �����/p$�����7/R�g����YlzAG�*�.qo�W�q�U��%�����{�6#�	S�.�G'��w�@�p�pA�0*���Ų�a�Z�p��]^GPOr���(Z������"MRALR�&>}<=����um���}%�]熣j�C��Wτ8��V�+��Q����QA������W˽,�,���c�%t�-����W�6�&P��|t×�]H9nm����_�ɢ����u1Gya�r��D�s%n��B��ܰ�f*Hc��vm��#���!����	�nG�j�����=�Ƒ�����G_�z?�;���D�Hp��zm��}�R ���~����۫�;抢	&��������dKO��U��_>�@��)K7)��?���,C��
�&�,�b���x.e��C<B6�Z*�m��(6���CS:�1�<L5p*�[����p(}5��4ah|���v�)c-�OKZTv#�5I�T��&�F�˞�+�(݃��}�%9��Re T����[Qm�\ h:�/��B`\" <���� 2��@]��z/X_8ل���rh�+얠���ΏJz=�Q9��A'
��,"�W��1OEGv����13mςV�4��*z�M�j;��	T`���Y����J>�1Į���m���ӕ�WgavjJ^<�^��p�㟱r���}l+bϛZ��悸A���n���	3L���]�3s�=��-��jF���Q��8���@��5����P�8\e�1N��x0m?�G��*"u?�riZ`0祟����[-��{fD����Ad/#��*}oۖ\�F$�BmÀ�rV�6eS��sNdĕx�9��:�ܻ�����Y��+H���m�+#=@��rIPB�;��w-�Zú��6Rp�0>��])\㝜�~��U$l&J��b��aA��&��3����ݔ࢞�X���نے&��u#�M>SpY��f����3��k�p�~��H�nG9����2�"��G)%!��{��p�g�<�L�)�#�C���a�!�#5B0�o��@���4��VR4�Qp��*'�7�Ժ�������œmq�:��&*���G~�?K�����������Y��ܗWDQ��4�o�Ip����{�FᆚyC�2 ��r��,�������H�d���|���A ?G�@2�u����V�Hb�Y��1X6)��֍� ����˞|_���b�5��
�[j�c�I:�
�-?�2*��Vj\~(Z� ���0��?��
gCA�u�8Siۇ��H/�`��T�j��u���l�����d�]{���+#t3�� �xe%eï�Պ���R�nNJD���C�~Y�˶����s-h:��q %�����|@�.?@�ʔ����$"�"ZAs�$T�.0��h8Y�h�m���-|P����'BY�uJ��~�zpO��P%l�.XD�c8Z?'@��O���	�r����6�<_A,�kJ �����8_�����F��B�6�#��]x��|6�Bz�b�o�X��D�̜��?�ҁ͊�X��w��Vm�A��,˚��A ?w���*d@�[�ﰭ�O|�W����^�9��u9��90:�R���ڨ�Wˣ鲋�<qd�� �wz����R|�K�Y�vF��s@��}�=�����aN�{Ne��j���y��E�J3��J[��rlqx���d�v}:�������Kf,�
�����e�ٝ~+����Ki|3�p�j	�TR���_�V`��."]V{|a�E�`~\p�R�jA��;��P}�/*�ոB�p<��o�W�h�2�s�G7���v�߸�m[�)O@&�����=舔���^9���E�$�`��䎨$��#{��~bJ�[�s惝V�w�����b�"���8�4.�Sy��<p����v�ݰ��K�=���n���c�E�I$��2� P"$5?�0���bxk=݀J-r�d~&T�g��QRO��ڀ����&�wQXmi.6�,��rF��<�����z���j�ec��ڊC���f��^�D�Ɛ&���'�w�*u��o�(3_��� �AY�eu��
�y.�2���i:sv��Ӥ(�dW���bxU���5	�3;6O��)_ꗅy$��P�s	�KJ5�Վ=���6�K|�/耬�|{7d۟t�>��[��gR�!C�)w���5���7;�����fŖ9��r-@�g��r�
'�e��fYqFH:�.^�&BT�eR�8�M� %E.���y�;��_��t��u�o���:��Ag�t=��nZ�f�خ� y��6c�XV��S���-X<T�b�V�h�8�m��������d����ߟH�nu7i��7�{��9�O����U���������V��x$D<�ܾ%�2j�J�_��;���V�v5���\�����q���=���N��N�G_���R�����E���o"�0��tV{�c� ��=?�9��;=�%�c�&&!�u����.��)M�.�#��̹��d�tj�"����Jw��m�(c��ɽ�^�3��m�U^S BpeA 8�b���a�5m����
wC)E��4<�jj�Y�lU�k�wr�K�*=M���h��/��P�����|M�����C���"�1�~���\'q��(n@��}9��:�����'-Ub`�P/B�r���.��3��d��_����\V/` ]P�j�� ��Y��#����!(��X��)�bˏ��5����Oȿ�x'��2�l�
G���!���x诹�	kvt�fC�I�E�Q�/G"��xj���\(E}D+
f� ��>^���J��J=]��_@n.hcי9����(�
�[�{s�1����UK�S�\��["&��z*�^��>��%Ppe�g�3c��q� �#�=;Eth�fu���K���V2�w\�*6KYaE�#CO�#M�D0�-�d��k�B�L�l��6l�eP,���"�F��$��<�&����z�h���x?��:�n'�$��s�-F-r@K���r[�[.ǠqQ�O��V����⺙��"�w=_&&�kz�jK>����<E-e�]+}����ӝ�g� ����Ȝ�`����G"��Ÿ����Gڡ>j�v5�ܰ�s�Fƞ/<4+��O%���C%��(�r$C��Sg�cC�V�m�ED�y�Z�����rP��,t���!{w�0���/�v�=#w�Ӻ-w{.�p�nNxX^�,�c�'_���΢Ե�$S�����߷�P��k�;�ꎻ��Bv