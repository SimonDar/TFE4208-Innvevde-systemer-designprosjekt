-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zl+jz592E3t0ryunoZpjG6IMV+EKf8C90FZgGlHsF3Bkxx/an2+remMd7b5KcqsDHR6wrg7A+h5z
4zO3rJ5blzpdkY3aJailvju+DEODFMwn6DH/DIDZB3RVchZo56B5LaELJ/OUAgwy+zXwQiDZ06Us
dx7oj8yu60DjDvXJhpqNfanB4dD5c34L2G7IU7/xi5mJSov3RabcdvlM4dFJsdaoV3K1ylOB10e5
MzA00yHxkGuHrLupDVkO3dVZwUYnlQUwtGpn0IONtCivbnlPukvEItieOPNHmVJg+ZvByZvuN6L1
iWG3f3vgOb6L6mzmT7fJ/xAuFBBPggMdc61UAQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
0XATlFi6DcHUHy2L67QHP2uTnq369b+pOgpDr3y8WDkh7DcbL1CouzUubTA55c4+6qduUf1qhdho
BpLKXxmpya0dvbtYlU3ocwqMmNkPn9DgvTlnBLAAACfmecRjS0fEZYUzZQn6WLE2JXPllJMrdXSV
ZVrttJ5ViTt/ao9BFl3WZ7Rf9tPPQjkS6GDXcYaD3JvN5LMcDJFIhXHUY671SXWwmcsTExocK8yD
T3YMRFrJTalXvKmcgStGddXNXOBEQUkXtmO5pmD5qXOh1Gy796G3XFbGmTJMYjrvWh9gW7u4DcYt
CmdnvmDTm2UIlZDO98hnTwZQe5p7XhAwM5O4qynUBmw9riF/qyvar9nFZl1rU1Vr9duD+AKMcP8o
LRSrricqmrUX4GvA1X+vrA6MQVfWKPcMRElKW527BXU/v6KqLWHQsuOYhStGurB+O2ojJAUdIsCk
azyAu4CNtya4AGJ3+8QNKW0dVQoyFgdIv1CcV/pDl9sRCGkbqRUh7I8+lAOyaHBZUQ94lvdE0q0i
m5vxrsH6N3PSZo3yx+hMsiRL/OuFg5sItIo/tektpl2quKk206q8TW3RgTY1doQk955qVEBNwF7I
u7NhSwU58Mru7PaITlcnA9u/aV2xVaHoG8wCs0FhFYIA8ZeRh8U0ssDsEMQA8xhcQJKVbVZeptTK
EPx79fOmRSk8+dOENsJ01EVjUJOBJdiL8QDVUtFehhuTK7FQdS2eAnpJ26JRQv18GivAU73Wu/51
GagOdN7nx24yUL5hRBrZo1y3WTBdx3dFOU3Ws5Fqc840eBvfMeegMv25kQ44b8RQbBcxins2RJHc
cA8LjLryPJat2r1XCmdUx/zsN0GCrC3V6Y85ZOz0NK2fU3FBYnf6RrleJhOgbGAYdQzbidGYX84N
rrh3jK4zMV45p2non3jR5E9MT15G2wX4laxM8E3zwqYOoWzd0/FjHm9pHLlr47MPOlXqC8s5vU5u
ON+YACQucS615M4kYhsOL8ZxY7YgxleKJM3PFGfpstiU3Kzvu8qpUMeyMr1sFkZoh5Mjl0zF1VBz
7XJ1QSrVEIMAO7M7pgVH9dcFf72OH4YCjwlZw0G3L+EtofaWYedu5+7eTClIvl1GDRTJEV7SFmO+
o82UDFJW18NRcjs0RKg/oKVhnBqr2ci7AUYVvFqF16lu/JOgAS8v7RvlDrD5ZJFYlI/KXyGXb2nL
nIYTUdWdPhuASMGoeT4latekXiIPf1hEBO94SbjsOY1LiPLFfz5Rh68zhHAHzQWffSZvW7GSxb09
qGAPFmKVwRUXpYs+I+YmBmZfEi98YSEMUMj37TVKQi0mO9VYGMJ1Ed3+V9i+qqOWmAxIMeHmzHwu
Vp62c2LuXUnsHRX9B9oYnFDSXHpRsz1no7fPwdiGS9EV69MoDbgBXvCijhZ8MY9oTkiXp5rvnenC
d4EQM+e3V8FD98M4tsNs1GUYET33h5hP5dzRtlBKIjiBiNAO1eYh764/Hm3rp03bopXRCS9q0iHm
Xd43l5Ak4yO+gsV7iKcS0DjgN+EgNhO8y8JL4rPfkBgDVqSwGJsIEfW8T+6O/8DEhD0F2HYFLK+5
91paz337SAiAc3oF+zK9CEfvxmlNMfNQpcXuOM38KjNDMBGV3KQsGbARg/qb6IExNhIOXXQfp4dy
4iqGpJAswypkKnqzKZXjiR6SDoG1wjXl5H/Bu8w9kqUo7wiRnsg5jZnnw2CV2Wf0L6LwVzhRurnH
61eU9mUlXno4ELuSLUDlBXdXqLpEQNHXkmicd8QbvRMVg3Bzgb+9QYHZ6R4E+jIfK/5gJCkzlJCi
i4jX7fRYisOyUd+/2SZZyIQIiMsaMbdwMssgDy3nuMvqNPx+vcoFkdr50Pr2zIS6atzjV4CK7BBp
kWg5fOmpZxv/vny1we6t6yGke6HLMf9WWixsuTjVMhl6JHBbKxB+ZzBpyFAEXQD0aTqSzMLInkVr
C4FSKfYL1rqLYn/CBb5mWr+BYoY82U3ltJgfhYNQyrUF2jIRzETARdvoUaAySOkFaRRGUZbe8zsT
lMG8AQ3fVReAvjCG9v0xMYQ7eNL4A0QGiwB57tvTB/59oEZYSp6+7a46ggalQAYUTOHyU5MPz8t2
md0HQyq0y+OnNt8E4CcInoTiH3/lBNZ38L5ZI9DWlSGbB1UPn4J/6WPUCawfkabw5Amr6Bcvg1BK
ARS9Fl291vBMzYz/dTu2T3ptX/7INiHv7cdGNwsNaK0d5IyDbpDsHF0Gjd/NuHqUnTy95+iHqJWv
Q6BKs/NuvMny/MdoufA2Bq9Z0KipqcmlE2yw23l0EynXYoXiSPZ8LY4bWWz2pDNVK2mmjv6J0DgK
VhRtqsOCy85XNRpjpd06/cncRAIHpoZBnUy8sW0ZPcRyRHx5iYMoqksbkQYOc97Jq0MUPsHasPz0
BSRoXk4NyaXquaJoBuI722l2kfFGxny6hS15+VhEKz9ZlHyIgVGUTme/mkH9JFVyGnurXyGoIgSz
gXCcm0++IK7507k8trZTPjwJ7yKsrINL3oFZbteP5ocrGLnma+kmJ69NOfJ5nZrTMOx48KUMpZSs
nvwJdAKnHjAb6AParoHEWfsJAZ6NzLRThR3ccGNJBh9Mupf5wvOiHZnQw3oS1UiUpbz6simtlGk1
T1iDqnsMrC9/iMXQyn0MJRp2nObNWAAx3/AIzK25Px0vdlCPqQ8dFaaXmv5C/9wB2MoElm1CtnCa
6WQqauPBseWEDodXRuBSF5lRXQ8mYiuJNaWeSIgnnnukhjD+OqJr5Co6f9pcQo3N4GLByFa628X7
n+rF/RqGrm/Nz8f4EFVvfVmef4boulqK+zMig9ynKsNxCpQEjfT+EseU/J3Bl39xbIzMKzvFwmUG
8VejJ0aWYqlLP1U4cxbI9Hy1E2FGLmcrM3Wp1JAB6oGo0sz1+KBuULofIE71FbLR5FLLVF1BSvVV
K308WPQGC9QXIAJpf5ZoUwTRo2Zxl52qyIiD8EBWPUfkqX9oajJ8dV314xv11L64OgKJmQvSrEWK
qJlfg398PWKdIFRSTQwHW2+b3j+oyw9NvdJUymCht65nenND+RRd9yoQO8TXGF1u5EpFkQPjpe6I
3f+NMNnxB4AbSPO55U+rnSxqGpHtdqQxx7Qm7V7GAkpEw94P1goOId3deNkkpFvm7V4lHt/w3ohV
z2Ft3Js6qRs8qClvDPDrh79veXR0XBVzpkrKXjPuf+KF8f+CdsRAnVCG2m3ApeqRdpFaP7HIDfWv
uSzkKSNmDQDV2Nqgx4WOC+lgfdwc87Pi41a8eVOHeENS893w6tj9srwYpLsXCZorDVd7HihT1W/h
ByfhBN/DQgQxdwBEFkmv5Dx+OfGbVVZkSC2yqUdG9cwU/ZvTjfdkhPzAGWrFIf1DVkuQilnbWCvR
wNpSBxwTyitGkWTzyZ9rr/udxnqh/8i1CCFvk+NS1xA3K+jFQNkZpZx0phWUhQY3FOqZpJ+XIcf3
S9U9oqhrJ6El3SA9DzrCOx6owfNQlVEO+fw5txsM4xPylo2czDvSVKasiS2U8dyEuMXCPre0CEL4
c1L4pUPfGU+DPF945fMd/yob9oytQOA6KdPhhLLGP+CrDgiUfXzknsTjOwPu8zC2d1VhpAbyVEPv
Jjjr5sL7cSFbrzDMVZEJ3/Ka6nlsxbnnsm70YzE7zK//tiJnr9+eVgMjlSJR9/S79dbj8NZCrrfg
aCZ/EHTQwjnGnwKxdRtJA/R5qWUvr31iXXD70IG+G4k/m4CzQqSU4TugD61K660xnmlTnsgABnP5
WyRPOHLaa89AvN6vyuwlZYsIhTl289+vl/HnEWHZ67Ua4crrzumL8FnYmo8r3i+HbvthkzPreIb4
iCHCden+FrASwpCLvzpxBz5Eoq85odBFTozOIy7aJwnWsPaAOemDSeRu/nRw1gPQZlFwKURnvGG8
y8jnMba0w1bqLKQnO7zKNI6iza7BuQq6NZ8lD+Fr/QjOHtWUHCZ6ue45Vy7DgR6DdPrmyncQs7hN
yhEZ0VhTvTPwoF6NpRaVRy/l3WZPZb3bIGqalGXd+CjjyHjJoms0Yxo5yV8ZV561vMrWo1NZO1yB
lk53ySE3GDrBJzS+n6bF6xqaLj9w2swjsW7o1aeNFlJ+R3UrPS/gDP4Ukc0FfjWJxktsIc7fN9wr
6PhoANxPcP4b+YBKn2fMW5UJyvkSRn52OE2W4sWtONSXJq7keyHkeuXkNivyIqSPvov6QP4pPi33
its9U69L3pQV9X10dUTcyhyRpD1xErZ6mvR56zHINOquVBBYkygbGWGnTS4dH6lX5jnKkWcf6Nr6
uike5j9bqsTj0oaS7nrmyxI97lSgWbfevTWhpZWY/FZge0CTj4G6uGS+qcW46jKK80/O/YizYFlx
/pN8j4eaE+ho5CQSD2WjoNZNKJESUebDF74ZTYNMGZeX4CXiGH0n4gt0QUQB6uSrSuzoJqg79awF
IwIQCmIHSu6Ob/nepJ4p/QP6JEU+QaHelWkW3/pn6vB+lLrSSJH1VHGvwEkU5ySw3rXWFuKeqG1U
/NG2xZy9Pb+e/rUL4bU6Al7+GPBNyCPS+g89Wdb4+HtJYXktennSbWhunGAnCaZtYjQsWNWfpv1E
ErF4TTirfpxJCdAB2SLnjgnYarWJqCxcHyIU3Yho9ee5vqvyPK7XbTFwdvtc4Wc4KLys+ay6aR3M
/a5MRHmBMBto2ErBRHFJNVHSRMhVRTkza3iEw1+rBUDq858iMHuCV1PIGeaV6D0DV2Yg6A8e+EIC
kE0fp09q0pb6BnrN2HiL1GhCysh9Mj76i8vcg1S8dukelcGhngR8DelM6orZALhf/NMykJNj4ykR
K9UYMSQzGIJ3dNDQmsAwBLDVSWBNOrCqiH1wPd2OJRiTrrnYcTxgABHtZII8EAmIclnbkL0wjvMC
mkqRLArKU00oN+iBUePk0eHdY4+RAbKyETlFaZQJX1oWHgcGbbnkukAItbKG9eDTAWBETtnywdbp
Lw7jYpmgGKNmeCz7juznuwZlW5SC/0CLuQ92qO/WFwtvY8Lg7NAgB+NT1OAf5NH6Efky35jsRYyy
HOgX2+H4K+utnZVfPFpm9NkuqksjEYiSGWVO386RZlpBY5O4cK72GNCoJ55cvc0WOSBicN8ZrjbZ
eoF/PwydM3Pl/tGr/d7Kyra+QnBseU/voUoeW+Xr8pBMfyiTF+L7J2SNq7meONmAkQHmn+9NzlYr
EeEq2Dgy0YF/qClX7/RDxfC8QzGUtiy1j7wNS0rMstfPm+NZTaRxmy3VsHOd3IE4UtN07Y/rNYB/
v2LUMSrHaoVNHzDqaXzO9RZChNnR/AGkAv/Dgeq504YJqHWl8KD2BYtgL2ntoOYAX2AVby5Tqe3k
lE/Go5JiuZ9dzL2P3R84MgPkDJCQL2r2VxI77sMMWCADsva12ON2LuovsTeeiSqqMX7fB9I4U1fl
Nr/RCcH2MOjm+QaQlZnglm6w4tejlkJC7UhgK+snppntlnj7H9czInSGmYrRorWtN9t0tx85Ul5E
IhS+ZjS+qI7+A12+sbR6XaP1My+3UolZxaQMwT6W6f/Myk0AnCl/jzCrmPAUJRAGplvREFbv76qc
nR8uw8G9PBQ/teocbFLkNehyDQ7GDHjUNwZg4vLsORdA+mUqoZm3fH19KtlDDbQ13Hd4xCHDLtwH
0MffBKEcfBwjYm5xOitKkzG6HQLihJLw229uRPiwsnwbxkrzQaWK9IgPMORQhVxqOH7oFGMRnFxf
pa7L5rDH9dXDgC1Mhvxtk/gFjookAlQFl+IH+bk1WF1Wrb45/q+BifJCwtl66+1Z7Qx41QafS7CA
3tE0Lnj0pbrIpKXj2eZeHbAZ95G5JFjP5Kcw7TpBTAYoFvlkftyNUApJztB+7FHTOPXV5rjFOHsj
CoUW31brCaoSlVHpbv9IpI68g6f1T9tdaYmq02FO6TLbCv6xLGAdA7bFaetlRc1yi7c+wRJLMyR/
m35igYK4eowWmZkfCjH2TPWW+vTXAyDV/+VFVxr5O/gJnDyIie1QMkGVYTfsh8c1xl7DQPcruiCD
hgJ1vg+W9/gjKANKlVXRd8Or4xao6roj+G5VERybWO/zc4sw+F8MXvJOc/zd5xo1cV2iQPYEXLbB
91FWabQ8wN3ZOHmow7YXDcUvQwsNkKAGcV+u4M/T2lhMXZRW6ftS2IH98SulswAlEkJdWYyE8hiZ
13khiFcY95b4OqEJcHiKbBFaLLsMPfHoOegjtyTs2hQnI3pFrQPiWEj0Am8RhnFUQJ9XfO+E/V5n
6qSRAIMkAnyYbzp9jFq12nq87PQWu/XkQbzfdJsvunvPt8XVWA2CwoUedjs/GuBDgEQu0Q0dKSHP
CQuie2zQ/H+OGsf9RA5MRZ4vQlC9v/zauyAeLbHlv1q6eT1oFH8S3CCVoa3r0Z2k0nzzgJL/sel+
et0RPJdlzrpOui3Dh2zWMvLl0wlaTFnpuyWK9k1OWTnv0iq61ZV7qoPctfzFE80btRhbMsXxxD25
6HHEU/LdhGyK5THUddIUlQ0GgUuNeM1i2HmUnKDEFzNbsJ1TPsG24HqQXBekkHIaKk4MKc138R0J
bCk85DQrLIBiH0kPPbqJ8hHOXTtYQVccBOWuM6kOSwXQl4FGQM6guApFC3JWbdRtQN6THCYyhEut
TYPUl6VbqFy6cTP3byrM/+6WdlucRLNWoUdb7caWRxQc0RCBVHZBITEb/OIsfJ4kIp0hnw1KwSoe
dqh3B9mJJXz2iRa8RIRjWcskreeC/1Qsb+pAFERVisalyue080nbjiGmN7tbKlYN5cIRq4LyPMnM
BepD5bygnDz/I/hjoPk+rddcKw9G3e3EWHSeNs1wYF5+lMLt2haRwLZjTYt07tK4/d6VRrNxfocE
KjNyz+Cl0scK9ED3AH/RvgNIlujjrIwtAaC2RcSXi3meuWn7WkiQlAM8xKkqi7veCcBrSeTLjPjG
HyBrIbZdTyRBjBVImecleGd3OlIoYieaNM4QHP2lWN3SIMJuW2934pQdEU6iAybMSLFlcDTyus16
rEjooKBgautUI69N9JE7phJPMzHptRjjUbnQZDNPfTmijYMr+93jWjbUIktohTwN1FgIpiWky0T8
camjouwwqGuWi1n+mhvUl4UKyYllcv6Lt+li9FmrQkHHbmBXxlR9ZfHGPNQMnaXnogpDJzZH5izx
fUS6bBX5iBajmPhPiukzxQ1VcM3OGaPkOApX3Fcg6D7E+g73HF3r8hQqoM1rzAj8iPkuYbNWVbMj
SJtjhSjs+pkOGlJAL6EPMElDDGbyfKoRduAPAmt2OzKgHHX56r5R5PkWOqHf33khuc7UJBnGIXAy
mFL+6T+gT64CYxulrIJ6VAF7xAjPHldhkBAlmw5DoCHsMrjN9+pgFhAX+9pwDL/h9eQiu4zlpcE0
AmtRT/8aeKD5Xyw7FRCPxXyaV+V3MVzlwhMDUYLtlnyDHOJ+UkMBJIC8HxLXaqdGTT5iTzCiJmgl
VW01qa0YCULSckKcUEiJbaPQau+NikmTp0YeQ1m625tFEcMtlBqtXKgryb+GFmbSIWYkDlX3j+ER
y/HV2EkcUMpn7CbWBTFNJAs9r6p0Gmk7KZBFvesVyCx6RwTeTvBxDLjZzjjliHGMhZ7FBijJhF7P
CtNEElZN7OTEsK0G8KDXo6sCjL4pVfDDTXAkfSD3oTKWXZ5FsYEreIxlL2Cdd1fN1aIIuWK1pYmE
Z0eEbykW8ZqUFrBlzqUX3g282OymMyI7/LQBq0vsDzl2t2+EnjnCIAiltUW0OrcjrHBOet9QCnkA
sGELAH3KY4XXfCoV5bNzHb8gvKOYo6j4rRNSWzng2dGfx8Q5pkrpyfEl0AD/pJN8/6lGPZr64AyO
epVQAQFpCBWBaIoR2Wpq4R0z5EwW/ZVfYFBSn15B4MXMjL2TyW185QIt2TZYOJ8bmSJiPHZbvl3E
COxSTpzZta04gDIh2wEdHzzzW5ZgRUgiM/YfyUUeC5jZmZgBgCs1CMu0PWrulgoW8Q1grDU12Oy9
Sv7l7lItVY1iOC+kJGIWuK2s2cvxFaW9Sj3tWwfJYqVjU2oNzRffVxjh23rN9J8w+xfAyBX+/+cJ
XLdXgm8H9QutyTSW6hTfbBzg5t+52O5iVd2uGfoBcCsrnKC+MvH8jHEyO+06chbw6/y5OWsqV34K
CpEC8HIItv2vTUdyfAQb8HhT9m+kiO5ZTYlEsSnQxitRI1QlxnCiHCLXgqIZlqr6dN5GgrPreMrI
d7agreDY1lFFRggvRsnu4r2rccoVrZHvsIP4LbisNdn365mcTgvnzFpDBq9LubniJkMgSrlIdT35
GKrN0Z/Bn5LxR1wYXuZvfkiBueyCChLv01bidt91A15LiwLx/hHXMKhmiQVHyYQrELcwoScju4VG
y3soyrnMIVZgpQXQFUleHR5NO1v4WSbQw++tw2PezKfMBNt6ulIMyhVwCrUxTkzJNfgmmyVEcwHY
wFQhrA+tfPM75ATRadINaEw3Q2QlvKAq4pdyHhsrfRbF7TI4ZT+LX8cwCx5qGFleEVPE6vX2ywT4
kNFOl5wDo7kK/RRlFu18LR0mPc7w8rSq35vQ/Ktoo7lsRM5yxBMhorC0svMIH/XzvN7hdOHGuvWg
ziiZg1wJt0fj+XT4vlb2OE6PcR4ysSBuroxIsCDgzizxnEzSI1m+VRJFWHVVb0FCvZh7q1BqjlPj
EAQBTWnpYUg1DGjSUkbL9Xajh1kjsUifvL4nLNxQ3IAXgO3t4j8sjk8WkGJSXeQxK91CAzmNzj4S
HxJ56FvJE1B2OsCKIEpQcvVeT73FM8apcAhSlpX32frOuJigOM7J1PFC44ZTxkX2m6yaDkcGAfH5
rv8eT0j19lP0PKzxROCC7U1bXTeNyit1rpC8NI5Sn8hPxSjovCMYFMWxTZIy1ceN9E3h0kuzm+9V
jFzSA6HcZNwnqV1yq3pG1OwXVlRgE3ybCUJGFAOxa0OeOQhyTwGQf8k/tjIoX1ZMfy6O2+EH8RKy
zIaEaAOpdP3RLARYGdRpeIurxjSiXBv230OSNH3VujsL/1egiCTrPn15oMYH9gY7bo6Yl4f5Coid
pw6dP0w0Phvl2kLlMn6Uhb7iqZiaDHypk4im/E6+0GTyzWNP8/OPUh6w4GkLNtVGmUsVndazfGTB
3wSjlwDMOJdNblKzaRa/Kgr4pWOXfeLliBHuZx+zHl92sUNCbOrtswhjqd1HsaT2dyU+Emr6K34X
vjnBTCfhJ0tjvTkXHKlBlN/4CcZyIxMEyvehEYks5JknIMsApz08LFNRdkoHykvTC9qBb3qmtbme
m589KwMwLZtzzNBy/hJcz822tUptW+KOEKC0dfAWWcHHITddg2ODtaJ2iHldK15N5k6LuUwD7CVU
aGQqHOtt22iX/jPyiAcUGAHBZOg2EzpMZE/5GDMEYsVbGVqsaUOK8Y9TENuysITqYZpcZ0jBFPoZ
Mr5fDaa3VY3i/sDYt0h/zjY8PAhkWqGYRllUN74uA65O6JWvPlMrSo3MEcVGORkvGEs/XmHYPDAh
PMGZXq8nNBjmvcg7HANowejpWtP+qX33fU8giXgbo2kwCYhsIEsECaIyYtyoC2gW+MOYVAU0hsUX
/6ZcZIo1lZCzc5t+75mZ0QzNUYKpC0BTXImkrKRIuo1kvdDUxnXxAoN/t5Eqcd/8mBxxQosv0BFf
KA8M9sGXMZxyiVDl02qrKe5p8Ur1uwnlrXnPt6gD5sU8FYjeLdxGzD0DjpR9MOZOtclzE1SGHtsf
gONVLyjCrfgy+YriyQPa1RtvvpRoJ/LM9T17QpUVPLkacBXIVfu2m3dBUU3+b5KZbjVkrQXff2eu
vLYnEnA7fagzEZCtYOT8a1eGf+8LWNzsRveFaIw0NLESYd7zNXS8smbfeUVcvwRaKPHM5rt+FqCd
8NNcmb1rf6tHxnfSGYcg4T2kwBGHvA9WiHgU/5XqCpG5RiYx1dKCJIearTs+FKHcBj3ZdQhzzk9I
NhVNN2+F2noy+66ki2ezV1q/iXDqV5eMj7GaOzefON1QQfuet9TB+Sc2+zy4Fai55fTItQY0yBcB
K0+tdiXUvQjjzbEfzDKtddm+fLSXyCCV1MZwbsRuIJjz55GxJQTonbgWqs4DgG8FMgFEso1oVRWV
M7qUJwMHoxqVfOCdY6QyVdD2QZwSotwIdVjjRPQJJxh/cs9MeXReQ+fJ+J/gW5oHtHNorIOCjO//
zs2+QhqumDtiaQYK6Ow6IO+Uu0JZ1VL9Vh2B3XasZNRvo+3WDtquSJ9zniTYKU4rPIE4GL7wouv+
IPqJQtvRClklfUQm9QabsA0sYOiR4k1MISluuK1M89MH64zYqGb6X/JOFOLqAk6geitwmSDkaCZN
UF7hO9SrQGaOjFlRVd37sCeWWgvg+U5LVGdX5b1kh6otSdFg0hf6I78FqqjaJvgEJyogSYff3n1l
R5qpJpcOjHILoEiWu3djsHpm8FtrBd566eCkdhIbh4mDzE7STi777eU6LBAdBVp4LYLYBiud/HqC
mgVNX1fjKyc9l2+l0myj1hZWSfg6KAuBKF9AE5oy3voKVffYMPOJMeL6so1qCEEaJzxgVcagEItx
XutCMxYi8RMGI+QMfiNdLu7sAvs20RQWSlVVt4vyU/ufWsWwqU/+jM25K0dlkDc1f2m7D3PEKNh7
Xql4X+JUsuAYCZHAUFnAopnkUrGSQl/gXrGyDynJm4RcHJiAobY7gHEdEpxJhR+FKQtgDr1N+S9S
IQyFihtFR0kpbv5R7vNmorPVqaPVu5PY4epiV519x3YJVmxLrOpTxtWyKnW7ixyHV3VoJHwiYRJt
EMtMhkylbtZbb83QAiqyOH4EqrMmx9a3QODuTm9wJezCARYesj82c5VAvov9y8ohtN4+RPK6q91A
6aasqf4cpM8bmYnhq1C4o3f2GNRJEUBY11tflDFc60D3Cpf8y2GSZMhQttCaJJhb+l/D7Mf7GE5D
3fLzw5owtnc67Cwz8D2XwZ9g41gG9HStEkwfruScHC+//4GI3v0T3mkRDrnsXfz0Aa9QNGSYkI98
rXZejTRUEXHkV55wKuFPKl8Ohb7aoMWlC+Y3L7N+Vyq+Z4UhHwMxwtOVavP0mllXi76pqwSi/JcW
Yd0BMB2JTuEXNg75FJH1k6wNb9r7OJbM8dztTC5DQS4eKpZMovezwa4ZtnRyJyzS78usKYGn8y3p
leUNAp9JhUtZzQzpZz/uLLo0fu175bX6aGdJLMNCq0uqFDzGMrbpRb5+k74zL3IC4bcLFK0QJHtX
BMx9kgdJiujT20/rpyQmpCOMSLMVISV+QhWyyTYTXTSBqlF2dKGyb5Tkp6Sjq2Y2huYvVj7Uvwkm
5vSOqNWD0JO0luLx60fF2NvixqttDRiupPF4GJGQnXZrXQxpzJ7tMt6jpTBTe3VxGh/ZvTjlYAoL
C7j1B02J8/8vh0AeumBJ2mNRPpHOBRJ9oHCjxckn9cAni3OWQ84IrwF4W4XhzIijlBTBX/4isduq
wEdU20oBMp3TJdBXbtqcBo9lPWBHwR1vj44/qdlW80B/RZE8Lu0c5kDXuREUEbThZJpTmHXXW8/u
qG8y3ojmjcenVx+XVFt2HJzTHYNmIGLtlA5KroXjPUCClIak0OlRgBes6skWHHz6TIDPa7/Jobx9
Wuk9rkJlrX8EKfrkuCGnsHWQBEMd4RTb2pv6Y+PEInTNtpQwpXTu8OmsWEf8nSlPo9eK66TDHauU
k7WFK81WFl+v/k58Mo/fPtMRss6Kw61XNDL2k3McM690Qm3oPdvpjo7UbcbuXsheovxefNh0dkVa
Vt25Vj1Rq/Jn8OPdGcEcpIDGbQnCFdVcloj7219IzcLsNpTENjKjbIQB7hqEmi6LOZtueEBDufc5
oih9IbUVMg8gBLvJC777Lv2CsyqKRH7QDeEdtirQoM7WrAznbmbwxRfAbaUqodx8bX/ud0rB+2cp
cm73n2EHQ1TfFW5ovm26DG62LUEkj2ZmgyATH4CW+la8jbPEOE7aCvEB8LP+q+A47m/LlUPtJIxm
9j1wUbh0GXUceyeC1jRT0tFixCXTZZYl1VlBTG7tdOjRcLT7Dnsxk3+JFPHuRnbHtE9UYS3THnGT
BS41gKtVFFvaW2Q1zrhgBEqyrFFp0F0ohXYubzjCTi3qAqWx6m3wCYvEbzAlqx4jfugr7nq1xDSk
q1DJ3Y8uKDq/rzoQZd92uR/In+VuUIgf6Rqdn8f3nVsKCw4WJK3n5UBhRS7vXrwp7PLuYrEmKKdi
If1lAMm9B8B5nG0RrrbjlYzPC458o6US6Y27iY/tr572yJQKSC7VxiConzdvEBUgxsufyDoaD8kA
tqtJN80zdWMuElqMhHKaQqi5N8SacbXPChNQrcbdQnYmNoyycMCoKpFVqDgQyMqP2r2Y/pr1mV4C
zmSEItcKbdBlKXFbEqfJvNuMzQUH2mD+1mdiQF2twqF9GRPuCzEdbtNe8Vt4jyfMoFJoD119W6Jw
RM1MIFkT/H9rxcfDuWk0FgkyCJyHQGjjkQcA9p/gnMzW94PTPtXNEEMsrF8vqAX3WAMS/JMHIWz5
RXdRztjbQ0p+kbTmJo/poZW1AeR3AshmyvK32CW0ruwJO0EVIzLFeRSo+gzE3sFCHu1+eh0K1kop
JsvWVhkYNRj1k7rWhLHSSgwhcHVXlURbQSkoinR2i18GI8p3ePqb0l8my42HllxgTDqivjhSH/Ym
KzAfh5GNaQIVebYM9T9HLKMliMS8rCF55FzFR5XmLJn1dww4/HrN0aqECojujeJzuf0WiGTVarrK
nJdj9YDW53m2gQe3JnfbyDvp0223Iy9qV9HrDUIVAnfwj32yaj48+UqgmjsuQsmcPbW4c8pUjiCE
TjpkmJ/T9b5OYKisjhfrIQLZ1zjBvqCtYLeFWBbMBYx1LbC5fYXYMTlb76xq4josQlLmtfuS0P4H
vn2pnWma2AvZGyenYk+2wFWLWtHVwKcbWV6pQUaCHMSv0Pdi+YE+vX6Tjf3L/sF0klUuPb7sfyOP
9Avezdy65XrMYJg4Q130+R7tmzXUE4pRRC+LbKaHYj1XZv1M/bPmFVFMAjIAxaXPjr73IspIXWEq
LMroAzoXiYByrv3lwq3ovEsMUPHlGWdFgEbuFD+mfF+n7itd0/4cbXXkImIikLReKsZbXICrlfCl
BAnZp0iZt/VrUn9HJBJFsfD1buacV8+lkN9ObZt2/2UhmLwFIiLI/z9H85CPeZVrfJdRVp21YyaB
i33LKtZBt6/Qco7Xh6vUfBO2zPO5lUkTddmVYxXJrvXuZG37Yuzur3nE0VEKIv46JMmL04GBpJi0
vR+/I3DBN4Fokw/qetbQoi3D4qSU9HyqLtdiUFx0MMNYuph2f5y+YWgGr1gS1LpYKLVBizk7bAP/
Jqw3NdPYuAdAGQ+1V2PcEaLdRX88OFB2rsQxAQYOI3tAzL5ySVQ4knDqcDDgywvnko1pGtn073sJ
Ga/X2Dh/t9NGY3ks+Y34mO/+P/UjkOPyJHIXkDo3mxRTD8ka/ohkFope323yD2HWfJT2UMZt8OeU
//a9zftCdABCp8vACRr3N0Fw+hpSsxndkaY10T8Pv0PuYhMJTE1wHuIeqIeXStD200ZxxnylADss
KySipJdXVVMnxKgCT4prbUbCMshmHXoPEo/t9+vF0rZFo8PwbbiQoZJZDkEFKhTm2YQCuF87EuR8
fHOmIfrPJXE7sJRO4SXwIb8P/k7rKUcFvKxe9BvJ2IDN3F0akiKOmtHPlTF7n8BfVGoYecoP3emh
YB7bfvLfMMvn+zxzpwx5WIpOX4gSoTCXSSZ1zHgVNlngKDZ8eQisqa7YDcuU4l0J/Kj8kH6aHMZ4
hPIJ4s8JharJUYvEMUtvGxQK8Df9D+r9UH0nyHq03IAWfmVfpW5mEitGN2RQXdpAYuMksDHKzAMg
xWIyfN1T45sAzlNY/aSfKnEbqj2VdNtzIClV0F784ztft8UzWMKVcGeJpp+G1mbz3/SHEY81jU1v
cMjRLXYmuUENBmpPTAYSqFlw97VuZtUdZIIt7/I58tphu6gc12oMPB1EObopJb8KJPm8O4fyB11+
fMLd6qJ5A3keV3yM/K//qbakbphgyNrQTy7XjKR8F4uWLRBlVrxtrbaBWJs5IYKUC9C9M4VLSCEC
5yTSsSg/BTN3yhVpGaRofZBZEmI6eSDOts3sTreB6KW40dvyH1baEJ/BDcZfUsahS3B4RKWQqoAq
kmnDXxJfqKBDl7CZMqHHkOdu5AFvAjKzSDiHg4CkYYsY/7Zd/GUuCFMhKSZT4v+qAdMnqd2LB/Kn
1El9eXlrTe1k1LeCHiN66LsIYsn+IX5cT0oz9gskKn4gYdwvPbLWj5PuQ4NFElLqoo284K+ULtt9
/mNjv+XDGb3chIzta7FijZfipnZOZ47+G5Vu9curgBBOAHpMqbBVVqUnnbOlpGT5EH3K1KixcIu9
6QF2K6nEPJcMZYNn+5eWtQagVtVHFBlhd9WWUmuk/giLp4hjLaQi07VLxIZHdlxM0ujJLn4rSkSI
rEc/iC3kOA01x6GhDgk8xws32DT8up3rn+of+EQhzLPKpHLK77CtAX5XDn1CeY+F/0bDg2CvNltC
OWmetetbqM90PARX4YNs7t6SftxldFUceHkOadkFgCrenK+FTV1MoWmOwWjIKAyCQcAo9u7KHhrk
prKz4gUCEJHYoWI8Kh8E0lg+A36tz3IAiyzm1uLLOa6AgLwCZ1yfnp8RPBeynHDBdoDf0Z+xybjD
pRLa9p4OnGPQmaJYqIU/NdjckVxfsFXlDB6SKilcY+P7FtMR2sQIjZwL43BkODWE8A37f9V9x1cQ
9mzOqp/ObaibK25i89nEDcIpQs4je3im16NTMnCLrb3zmqpCZVEclJhShd6bocScThyMnwKdkEzT
TTYd/j3SdurK44jlYTU6q72yYzpY069Ofb/jhy6B1oM1PJLCGcWqKFkSWQdxMiZMEcxqDDWJpugd
me7lkwVRa0Vmw21Kk9LrbbDd/BLg1Jzq8p+qf/NG6i7UeuB2nfF0iPh/P6TMrIGBiCy0uPzDtAD2
BORA9iLDS5Rs64WWr3FzM0JSmL+wfEBI/aMHUhyiL+MCgRa+wg/7s25nZS8ddFpCqF7Y/u/T6CRV
wXIEe220HFtvLoc7ez2ECR6jElR8LlsZelCy3rHNagSZZXGoIiOPKSaLveAkSVimST3Na5NaWPZ0
wxG30561nE6Ufpe3sUJUFcrIJVvEuu9kBQHGOqSLyk+eR4zOTTzoQFpBH0bHgV1fnGoug5NO5yja
w17rHzVAvrMMJ3aJu1Zh12f5N97CU791T/fG3TlJ+USTqVYDs3Xb+zdp47FnkLz7X0fcRyOrwfsW
4dTKXyfl8inSgfMjElF4tpJyFaZOl41wjbHWmoJHmSiFbimyilhzXKcLIa2kdWvc1qA7DTIhf8Bz
Lc/9jGK0I3CFvy7fVRJra4ryctwiTXVqOIcFm+Y68QvhbziJWoJxpUXDcp+ONZI8J5M79ahJj7H1
10YYA/6xj6OG4nVoPQsscLVStrncorbqgTixrL2vODsehX49HBdPiHT74smsCiim27zv6Y/GTIvW
zVq1CJXaUQj91s1B+asCTXsN1Q0V3L0RGBXXvVMR8R/YnmTkRNVb35m8HXtsknIN5aQz3DKXIJlM
pGjVS5ORqwLqLKKqUO9OGc5qiVYm0zcZ0weEupYNpZd65e9sUrWn0TjdcKpfI/UE0cZvV4oDmGr9
2TZ+3oCE7Y76zOvMa1ohr8mBI5UOosaExTB/Y+Gmx3ijGCoLXCe7D/dtKROSONbH+PwPWuiN0Qx5
7v6vN9oPKtPj4q85zhPA4K2X6xGgsaKCRLdR31OkZ3o1Rk6ut0woKPSfj9Ssb2hqCbNLafPJ7333
SAYncnRd8CD1HL3BSsSf+ubUdaZw3ZwCUMz9uthIKvnu65joqXoppOYjKnEwzMfytojnzRZHy6kh
eKt41xXbK9BXqWWB87i7h/Jzzy2csZRfNQ6ZR5wZezHEoPUpbU8DFdBIxPbChYW+oGJLHsjtcYYi
xaFc4qpUabDej+yLV2TPYmmI2xNZZPz7uLdTLDEhxuD0JWBsLA1XHaes0o7R1MJKerCOptETHsQw
WLroPFS9ENmZgKO1ptuRuGTTC9Db0rEZZ9dGtVFGEwaMxmjX0x7ej5tOl2IQlZRcqq5EoogkyEgQ
YzUliUozwDbNQRQO6vNVAn7JiKr+y/Ygpkz00zZU5HrGBgFiSUqRuNATAaNYfYYnx1aoCDUwVC1X
YLS+QTwcPMrT0rCW0LMLPYVWAtY6+VUNPrv3+oby/GicjOw5xnimfnPGKF5c2Hca7EmcQdp6dJQP
/nFLyJc7duLBFTubDIwYfjUEVPN6w1pNTGF34/fOYSDNlNoohNqozT/36aUuPrD8eTAMpFmeFycQ
cx62n5Mw1Pv3Xfq5kuTZs8GtOaPYANU2qdmH3EQsfD0OWxaSePahgvU3sAAh9M4P2TDDV+OQDP6V
Br99AuVkINpvN57anKn8BoVnbrtgb7HGYeYoOrJRNO3rip+TgbHUioZGj0RakVeZTp70stegv9ZX
M7MvOI9kX+be/FtV60ALBd9lSGu5Juoy9z0OMjFb/GiHHjxppZnfYY1sVPGT2xdQpXF57IdHEXrY
xwu+NVCJBNX7ReZsxTF/kw+fd6DopzUvvsnOnudKqED0kwpM2sY1IBW05Sz4bpKB4gWlRu+B1mBC
XX4fDuIXWAsJzcwnfhFiazS5UZQeuMNUNLEkFvV0SWt6vRo4ssDSeam15xHJtT9e3/FEVoAiHQ1V
pQo5L9vm4Lv+GjmXmXS6aNBfkYhSINRm3d7m2j/+csjQvMJStCo6y30PCh+ZCPoznWQTpqOG+E3d
507S1mfUsAOw94nOIWquralk1/wC5GB5zo8OHwe78hD7riL9Pvbh/uzxYBXF8wQm80ty663wG4Mh
ZH6BAwFdQ8qfjWWkezsu8eqzncmxiYPMmNA9gg8Tu8sDDqneuyA1aK4Cg9+dCbjV3h2Hs7kGH0lH
Xtu+ITFT2yX3mhayFmxqWis8iQz25YSrecqZ/Dk6svNWeWvetSeP3z52sPQxvk17R13+401ZkvsV
2FVdfwGot17fzjju7x98KIbFBZyCvDh0byXYM48/DmqEV3xSG8F2xJsKatNLP8InujlRvWIW9lJV
qZy8YrvMDDhPj+mQSKNVAkZwKTBZ4/Y8JXVpvab2s1IXug9mMR1xDXq/6ZXgFhevxlYbCQxtQjrF
1bv4rFK7EB1auIoa6j6T7y5KpwfjA8aakWyRUOj2CE8TIyTpkReqn2whn4qztk/aHNwJrQXPEQCb
qDMhC9979672enmR/IpyuAW3W/qmLweaPIQ6rxOqqoY105K8eJxunRs22W9H7h23SgkNiLxfTOBS
qZORm18LX6l4RXDyEfVvw9M+FdrKsSW/22gS1L5LaeZMQGpYrAmQwddQUT9mqDO+px3OFXHXHJEz
KCbloxlL4jKC6RDuGqwCZkN6OomkbDpfg2J/RVgz8MQUbsHXbBT9M5LCRfAGP2cbwvlLW8RZ7mVS
M0Po8WGTS39YROGu+wx18a/iyffO7OXequ496xjd0LgcfFYuhinWokOik9YBFY4UjcCGHRkenPaW
0LnH7hJ+LC3LsiRk2RXW2MsWnh7V1eOYknt+sCmB8BaqU1qQD9nKNKxYLfpyzeM8HepV26UNTumV
QT8Umn3n1jGwrVMkpvmy2Hg6LnwYMBKjPFgeOTo8Mhqf8Am2QzbNzsmePhUwBUgOs2j3WDWo0jji
Uuc/xyZZvpzpFHPLom9MDhY+MFUtbw8kfYmUJMv2QRcjp6ktl0Fi7UL7xZmdflknplalLUvykNCV
W4589w==
`protect end_protected
