-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Aj+EIck4hFtfhuFggliBM89ncT6YZ28JC7aVZqxrliM8/Lyr1RREyHBSqtUwQTpG/6BdM+tI4Lew
FJeJ7t3Zu9frtsdlP6bbD5fPM4yGrw83dv3nlqAmi6kM1N4Y7dQcwHSx+HTQBtqnMJxOY/gWvjhL
cs6n4WI4WhjMIRpjEqOeFa6xHy8Qofp8jZotNliJtCfYobYPHE75fRzG0XiEbN4ivKi5NHtjDLjG
G1gmTlzJ+u4koFLehACoRCEmB8W4pNRIdc700IoWlgbVSKUEILexwHdjVpPHg6m1QrFzhMA1PPF3
Q7IpHP+lzG9TxzstqNNblJVAZmcS2sgN/tiOTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
EnFToG7HlottwRXBULHKq8Qo0a5R9Pcbu9rCWXmRzAneiYoroKKNnryWYAY5ygmoXuCipBylIKzX
N81PS7T3WWzOOraYr9B159Pt0MdwKIDTCwIZ07hGASLzCJteQhpuq2gXZgAvQKI9R2PyCStJ+61V
6WiyWIftTz1qzXQ0xdrzcbqx1REfUlPkzg0H9EUO8eTim4dMFdI8EyQdNgbZXtpZd6pm2o49fFBA
njUWAEsTEssNudgSIJCy6xaRuFyVZJPLusEbgVZ6IxZdJIOP5eknfx1uc2YZNMUUg0nL5XBxDeRg
Gul4ccyVg6qaCr8RjzZgmRESOUcbQbP/D2Gd88UyMPsja+nEExbNg1fnCOi6IcJWLUxbPT+HJzxb
f7xYkEX9S84YgwRxvl3JDmEPrwIOy485fOanTIFXelOrhUUwGf067zB3rsziDxyYMdfmAkuqcznr
+2MTQ5FknqPAC2MpJXyLT20IGAI/X18a7+ZOeIyK9mMgw+gMqxafJYC2+6/H8K5F5NIW6+ZaMSV0
5jpO0+Fyx4/WeKNPMS1xQ+UTJ6WQTZGUeAjKef0shGqDcB75FgsoGNRIQOOOAGFAlIYISjsqMMak
TPwSzqFDcP9AAdwTX63W4OGMyX6p89TWHYFzuaYLYY7a0fCrG6y58ATn9rKg7s40KA/ApO82lQsl
7jfoz+Ao6u9KjGg2Hk+t3MEl4+uFPveoks6dg4iX7P7p3Mc8vUJR+/DJgIO7CrrLMeLSHm9XgO2R
drBFTYf5fRKV0m9a6j6K6ZWcciHYat0biXzWU5G+TCBMAClehHWrM4beN2REnUTE8F0ANmOusxjf
0ndEeyvDcfJC3X+Gcdr5PRhT7LVPJQ9KnBN0MfAWwWY+b324aRQIliEAT+HEtjEi+o4wM0tkPwVh
NrJIVDSWBP2730lGjYT8fVAis8+bqwKMselu3r+KbJiWYGfAzmffber+7l5HaAFEFjFOxCOl+XbT
ePsUwfekVzeNDpJP+wqpIPce3CYDoM2QIiN2z4sLkqJJIcDeraWo7MhqQc0ZqXo104teiNQ6enfF
wJ9DYVDtRPOiw9j8VEHI6pgxR2eR2FuoemELP+gFESYtit7Tw81+OMBDeaonnz8/L49j4LJGvWPO
SzIB5oO0I6pxt2V8RqAaqnc1ogo3T4oEc2GZ8pch1iglKxwAfBchvt/b9KqZTk7UuEPfqm5SVDtR
EhH0siSGerEmCi+KIEYFZLJydDE8qOKOEvYqHB1z4ROgP2Kn1SFJbtr2/kDS9wkrJaLqdvsHNF8x
pPI5auuHMvKHq9HL085OetgvVOuJXusGwY67xiJkCq9hqZ+N/Ys1wfvijc/7kOrgjt2D/L/+fDi8
wcBwHrFSFTnorDppHr67HGGjIFIjyyymgytV0ZsUQ621eYN+DJf4JhuG9smpKJY+gaHFTSeNpjFA
/FveXrVt2IONJGt9qd6naMCa4LivWkHW0UpOpBzyDndfV//rlHqOU7Ohw48im2XHqIXKDO1QZKYA
xngziJWGs0pj4hM1CQNk2QBTKze+Wl1kRyw6Bs0F906huxSto0HaAnk7+8wDeugj8+LqJJ7stHn+
EHG21rA/7KKjDbhmgI5PI6nmU9p43os0RJ+bewhdmoI0Bqrep9aPdxnWuO5m+TomVqT0f59mnpTu
l3SodIdsW49P4Hy1FvfXsgHwDV3IKswaIUEn2p7GvSXlN1VhP9ExkCQPlstiHfuJRbG/ZfuBXvxT
nDn53gDsERik+xjiErC9rH2G5ZM3CpBgtYK9UAWmjERsV48UXQ0/hP+cHpYkDFGG5FP5HiKOmGvA
KvsuwqboPVkAKNN582P3DYtmu3mmqcuUbDd9Jh9Q7lXhyZQtaGv7g54hSIrrFu8qIUgA4L1Jq6ue
7gdEpKz11LJMQjKwy1OEH+lKJgdyEaARfxjSE6mCGkFLQBDHgP90gzwBtz5ZA4iwpJtFtXSuTOCx
1lVSnHCz6UrGxRcDqzBVvLuSpnJ2HsmNKQgEAAMdHFJgkY8QNJzEutSbFFMkbJ9meSaIxVw/Mri3
WIshh8Kkwxfg2po1jVCH2N/QiIDMyhbqj+g7KA8XeXXCOAuDhKLSZC/OLvMDiOWM3sYUwXjeWMb/
bAPtIH0pVRABUru9S5fEp6FisbihSGsCpzOt+1oiIJxWjCzljqaaOvlzge1EYoyyaQjtpt/pOWI7
NHmMlZ4UzVoSu0HVSMLVGbbS37uGbDT2ZI1yOQK3geDc4Wr9vJnHhPDbKySm7TtjnYrmSq4v6Wf5
LmKZYSy5jQYounSBZ5A6wriPFsjZhQP2JtxfqoGjbn7x2mAS0chEuMEWmBOJkU401JKp854Wtjb1
UloAB/c+l9E3mAlESHlU0DMDONllAybZ3bp9HaC5bYquXcMlOFNQkabSzeq23p1nJG682TMbPQ0R
KeDYaXaQ51rigPxuyms2oY3TjCm0H0S8E6aX1IH0TwCe7QQhVx9FqiM80SJ7DeIAGB7eASVesoJ2
go6hLrmpne86N1wbJNNFD8t7qeJP4UjcoiPYY6ktarOl2XKKxIThHetVWcTO0r8xhzqzp14XvLrD
7nFcKCKal9dBVw26O/ppy6gCtCHLuCKLr1QcTZwjyc89nOJA9pg5EcsJqboMVbqWUpYdyWasqBKA
J4sMmSkNfWcHhqOUqgVMxS6ShAwo/m7NgL3bU/EDqg78qHjVjAdzq/UXD6z9gHZ5JSV1y+tzwl6c
NEWlY20DrqEVcRL/LYQKbrK4KA9aC/87TIMqjVO3/chst4Df8KyOzZagilxBDUnMEzF5hUQlVJI1
YsxaYD20bnHXoZFGqNcfD3+pCj4mHs4UK4zcgFpH/9VizzgbvxQ0azOrKM6A4C1Dn18LvsdIywxj
RTKW4gcMnZRLPWZUsgHLp5t5V2f9q/+Jl+fP3JT39Tqq9Yop0vyrdLcd3BbnE141aYx+92TPfuxW
NXE6RuDXSR9D0aYisscwR18OBUMC2mDWGoh+pZfz6I9qDgnYmYkk6GaTocCC963Pwxji4qu6Xlf4
KhXWZnIl82bIMsyFc/NqvDkMn9SGREjvEEk4Z5+Ux/CYWd7GBBtWgN5eHMg48SOiKe1BPG/boDCX
kVSkyhAQTzcG9hlqwjW2pJWH4dL7bBt2ZF0OCQfE2T2kaSi79J8j36Rs0ofzJzc0LQrQxJB7TTLi
JHzxVCOwkVMuLR7kISOLa4w4QKRSo4MyOSDSyQRSYq9ZgclDHn+MoeTNnvOV7GSkYwHKwOtfOXrB
AxCwEdnb/WnLd+KIyvcp8cw2agdM77KzUDOPnAqWXV7lQz+rHDqoMeTf8rObx8GmTzGQVAXhP01N
8RY1yUwmpw45xDxM2x0wctexz8+Ce/n/gmTa5J06R3hpghX2TTvDwABFRhWl7+x3AMgXVa38cHmY
cfnluYQEv8Lu+IDZpgCPRrM2Ku5p2LMGm9HiOkkBY15xgQcuQRHtGs/xM1ZSaJD9RivlnUI4fIB6
IO21+/O9689/99F/21jDgaFTz8Nrfnx7wphuNPy885szCDqdYfbjWwk5/xKf4Gp+LLT+/l50KVsb
wY4TceCoqXLWhACxwA7r2UqLleeFS2tswNG9k0iG7Jbmmp5Za09Oq87PsoKzniIQW6yesLVWgWpO
hMD2Mnj//JBAcQ/msp2NifRxjnzg18Aa7nQicoZNNbBe8vGkeqD0u67H5p3q4yN/upCiRc2ld+ay
30JcG1Y/9R/iak5qXN/gGttz4SN5SvbJ9vMR6TtnX0LmK8hONJifqDiqvGSS9a74mG0i/uYxNncE
+ogTJQZGomnuHP1xModS0PsTFxSxINApiib3n0Rk8wVWc1PDqoVRfi+S62PUS+m6Y0KmZ1bwBqjg
Dnf2GHrSuKSAwsVepqsa+OGIY1R2xFcdSuKkgTHpyCdXUYRDFpQ+O9x++lcrr3LZcRrvihrOyP6l
OcXuyLaYxCYXS6+o1bphuh7FWYWHREgNYsNsO4/cmn5Tf9q8f7U3iRH/4sHqSx1k7UC5aOc1mgrC
wPMuznrvwp9qeU3AeJodIHKU1EPrkE81qf8zg2k4SN0htLkTXGrcJ7d7Umz5FkDMuLmq2vbJ8mxq
WPu4HO69H8+ERG1uiR4pXpT/2iDUNKxjmAeLTVgSLokKIllnJPMB5si6/wbLwajEzyETnfTc8R4W
uCC3Dak5uM/ZCS05HUHPzy5b/Q78AvuDBK3kYlusvcxXH9VMencgFF6b7sdCGa7b4lNvlyV92btu
Vm5VjCosBKhePS/WBFm8HNtYfBGRG64tRYOK7pdMxviAoMvisNbKXJ4l/GKYHKsKXFFeH+J9inct
Dyura4j8nCDgwf5d86GRrHfK/pRX+thoMCOCM49f1CpFhX7s2DYuMJealtX8v3pL+s9txm2bzjPv
7x0kM9UIOOViIYu1mA1xqECW9MNNWXWJjvIKTAdGs8Fu6MHQF2RuePesWIAVG2p2hM3r91K1ePhe
T0IUkg0fMATmFkOI/ISRDzYWjsKdGeYV+hOSKoY6swjRDW8NZtbS/IkL2+/8bKaRC8NOgOv9FUR+
mKQC2b7cnzJKwl5901DHTLaZUrCHxx12pVv3MiQ3uyVZ0Cv8mP9nV5HtwjA8tYpg2aMbzaUDNes0
hB8R6WU3aJi5x0P9IbnpBFlxjmlTGuNilrUOdwYbTLvKz5KTaO5tDLgzFuOgja2AJxHi4soksPUV
nw5i42pdAjFBPb6EmIjb+McxaO4zsTHY+GO2xYuzaiLjalpXRq6cii5COX6PhEFZWdA8aQpeuYHZ
x6W2Y1jFGs9cwYZDNyImtgEZYlcV9XDDotJIcD1HrJCjT0R+BIiUgwwVY8hD0J9kc3lbAAnojgx8
/AmDWbJnE7wloKN/MycGF7LzqEVoq0ZCMHi/gkEqoMZvoeQC27syw04LMejd1//5YacJVruSjL+7
WsrMK0q7+2j1uB6ExdLeseXCsWKdXybncspwlwUmWwmjPJUGA+D18b8iS0HRs/LAzOyPYkEnLW25
l37MvVZPXBcnDBj0LzldtfyAG+c55Rkya+bEJFsdJqAn27DOERGQPXm5iPmTYZRbOakOLrL1n8VL
8rELF45PRErM6OJPMj1OTnSPeCygihMVZQOf7ruJmMXdbh4HDH5brg5ceUCG1td1y9riXOTfyJGO
fxsIShfpMrRyt+RJ5JTl15hJIfO/ioeFdXdk8y2lKVNuT7pfISng9waQYF/mcNKoSfVH7vaIcMm2
cDZqhCVDpdLO5G2SXLdq1WJbcZHtYWOYCgdrzsUi83FVU7HLQzuwLe8UUbbm8k2m5yrCxe5bF/WY
MJCM2J2Ekh+NIui+dWq7l0USp8V33PYLgdU2qkFTTvB37auo4WL++H8AEaRMmPXWuHD7eMbhbatV
lpL0QJsr+X2puzq/68ejdSFvTOb69tFis0TjDi9DB/zO6RX+BbSQMjvCFcqy60nuzS25G9wDjGQV
Q6pqCLvDWKZLGn9J49l37yYb+niStdFjJplx8GleiaNDYoKU/KLr3+Zb+I5D/ubBusCfd6u9jR2v
7rqVxaoS+c5lJE4PX459BpLgjWS2poxxMwCi5n2/5b8ezmsPcAAR+opp+1AJXp1U6UEJtf2hKOVw
cwqf/5cDSKv0OhX/rPEPruJVEjFyUg5kK5ZHk950jMB/5KabKLEqMC3vKsse23s2hSP3qRa+OvD+
GG0tCMO3mtwqHnDSdFM+NpYfS1t4mk1ZXVZBtyvTUq4oTvvoOJO2mrun2mvxPuNX9NRDkQjngjaY
V+japWk4teXn6dnAC9C6CyLfSUEIAJgG0Lg/GckdPYHcd+pNb/+gLUNa8uLHH2JkIQ9mva5o+e+Q
09uIDNZPh3oW3PQZBI1McFm16wbwGvafUXW795FKB0OtWLDJwzhd6h/kiOURMsmw+5Mde4C4kch1
Pi23t2pWX3YOr9ZKu4qbfCK1wADk8tHldcx/Elidr8QMcZtAJ5hdsl00e8gQ25rmgqduAh39s93T
099vfy+3fC7T4seXCTtjShKTLkmlpjGiHZgI6nUobhKK8weG6lRhB0qU29nPzUFIOU4hJsWhGJxx
GkPxBRVOtKVNCX5J0Oe3D7cl8SS17YX6V5hzL0sDpQtpIv4r7/HZhaYdyWDqMmDgfDTdyLqG/7qI
GLu/VekCHHPGTEZ9ThSZqvKdcaP311RjCej9h8Z7aOzSsHPA70icI8G+VrRG5AXv/2vwi0jRdQOS
AVLZDEQWm83KSSFVfTjgwrlnmM8Pf9iAO2q6xy6SDZZcXg5hPZoOV5IBxAlCM3AlCyc03Pd19O9/
xfTCtHBA95dR6beu4n4TTBkiZnnxqhkDYLE06ySuJsBTEedfwhz2DVIcRy6qp9BdJqjPU/uFdb80
bg1DIe4FpIbldsiLuXsAijE98JpKh4RvGUn68Ov6NAkRVPtl6fkOapB67u0/4QfW6B6lkr8F6K8x
1nA9B3Uf10XnYcVg2VtKnWc5kg2642Vc1DjpYpmdenWVq/hd2T8z103exE1LEJh2fU/9/2PhYZtH
dpJDP2lYzPickiYhnQ4lGq8BWSZ1Cc95EdYttwgXEztbKZxSKzPUCwEVWCCkfSdvYkl8OglKlyyE
R2pW3dwsOe/LRuizRhLG/pEqljQeHjsoE0E7JAblbd5OcQ5W8S6Sh3S6TO9Hh6DHt9jtrcNCs9s5
S3koAnoubjKYLbeqgkdkBnjzDJO80HwlNY1KM/dhzBy5UR7IupOm+0VmE1ekhLDk1XC+iEfvFtsa
46+va15roaIVgyI3BBwfp8go8Q3un0OLRwKx081s0QsZUMNs3zqx1ef1ecCsh2NHpGztqk6e1QfN
vxe7VoLlFt0j9r6hAj811wheWr626SxZwg4gMpAZ9y0FbhFMXBeLhvck7d3txMlxoN9hxBaDUpbw
F1LFnY+BU+5usJ7Do4OGvulGeqZeglWz7wS932m3zX+CciesVk8N0cHpRlvXEL0BG9SGMAFvL0lE
F1H551tevBf6HVjiLBMtLX3bPFt/jSmaCsMC60rFI43CJ+myLRq6LA/4o55c0GnwyCoJXzbSYPaZ
nMYT0ELY9QQf6UkUFFolcbsBJLvdkxsyP4Uhb3TRPNB82Fhi7BhjUTCq0V33hHutkb/nSZot8HDk
qpt2boSzmR88wYXEL+WuPfRjGs0rv5oIKNn/fNFeThKdX8AzHvwJnGlgppAA3kePGdomtmjixwjv
L7bzlwbN2EFAkZjlxyGicPF6CJLyRYPyNsDuyuYoIBFmXilFK8ZOHMWQITVuYNA7+Rk1FfrpyEyR
x0ISaxxP8mC7C1daA4+TKlCZmaVkHL6ITwdUYnzqPl2gq+mmBE+gMthwNXxmBRXePbm5y0WHmmJd
gviHn16tnCkGj6HKSYndYB1nKF+fPashOBFcJszS7YGHp6cCPB5l8V7LIY4tGI9GZ0zHtiRz/Zyi
uv95/RjdzQle5vo3dHOewA8/Z5/+++MUTR3lFGHaTLW6Y0kENQIQp2ZCiTuq65TrPUUQlvAsd0pu
dn0Jqz3NqOibtiJ67+eo9VJIrQArqIlVJMR4jYQjyNJMQwyVfYpTs2F9l6rOZgq5tXzTPz6wm1mQ
PwUG6FqFOdgB/rN82c+rw63djnBxXLjKQp74kxJN0zD9yn6FtCSEmJaV5WVjLCKdvbByX6f5x0Ia
shyhe4cnwCVTtPe4uufc5LqpKteOgdpz6yJKW7q+pO6PEm6pLFB4BUAIjSy4EvBHsyn7wkcyaK17
e4hZb0JcwuJjk6Po3xjmbISniejhvbTpg3C0OTi4GhAIe68IG0QP+o4pl4DtMQZhErC0DNGGESEF
5NSRKhB21dlthNweMw0h8LJ0AuXSEW/MZzeutgRyP/H0NTx7w4DMp9/hAbyXvabrXnQeIw9gDlRJ
XRcslsAv73a7bKGKWNKo3R1k6c53wk5cT9ju0NOM9hfbHG+Saf9Mvpgh9Fcl+WflFDG2V1omrEAM
3ViE22ZHkSVAPfYr770hEdJA+dpilmV+V5rvk8eKp3eQuv2mCmn6HNHBR8sjsWN+5bN7EQ9tKSSG
vfn0N6gdAkw59xz/GO7HD2uo6PdY1MpFr+/H5M0563sarfNtxeE1wxrgIAYNS+4btZjNzMgkXyuR
E68B3w0wfOrZpQjYKMVmCY1FI1bu106DrfnsAkOMhYRYRXj5V/qcjQOECDSIKvUIj+XoEnP4WpC5
lgyk+q6kSjAgyq+HiZO+aZRT9xhUXTyOzt40WmfWcsW9uB8KSMSUgmO8rMocK0CeiNuMExpS0Idh
yQ/Qo96kSQVq2af5re+yWT9jYrhEflQ8CmON4VqDW8nJmRruNzy4ef5va8caQJHOopKD3ER4qWvz
TJYgZY9PBPSYMUcEQ2P4J3U7ONSWdZtRXvk2kJPEth/iKeGmYYzUB1G2cEy/uoZ2HAAmfRLSbTvV
iddeWSbi9DY9ZmUzm+s3NXnc4jBkdyALWGDiEcFQME8+Wk42go+FsaMuy6E3B5qgnvDROjYQNnsu
97TKbDnqCrokca2am7mO8J6gTq358/019B3YpvskBiYozPpspK3ZlAJimE834M0wEzUP2fFFeXFE
P6ivicmI8fYX8NckxkLsBPrV4QOhNASjuGh+jfhFOzRODN9zgeFOCt8FnhCdyi+QLtygQdaO3jQV
7HbVVsB3xPm4zMz0vEBcv+9Rqxhlc/mkcgyYhpnIBIr0G7ZjkYVVlHmlasxKAS3PaN5Vq61z9kMe
8YLsexMlarqs6YcHruM8cBygvBL7ozWTH5kzW0DDFBK2llvQSesRT1pCaF/cpYXqF5hDRqJ6lC0c
mu/0ZuHcRd+4lnGld6aKkuvrsvNrKh7/WxQ+lD7UXs3RjrAlQfvcLUF5J18fcnWXXNWhZ1yDI3eT
K0ySI6deazD5OKW4Musza4QCbYB2VnyQupREReoaas3vNXYenqYuG8taPo7QCO7AQ4gBkVh6u58C
IMAnIzf/blIATpFzNBaSgGd31WNJJzEf2Ff/+DD/tVFyx0H+vkhecaO7VqLUXMYvnHGtjGhaTIr2
fh/wxQNt22Ky4EAKp7CYD/t3WcycI+8YR+3xjVQ2xct246uCDTSiHvYRBirsddPTQh5KZVSBjdWb
bagfKYKGWXtZwNaWjYq/QOecJqbNYF7q6oX39bSjPFQDJw676uyA7nFM8xIpbc8lgiKfAKkTxe6Y
VVg+PTGeXkQ3rZAPg/NkW3JpdBpPZFrp5CSPs3OX0ssJ1gCzdQeTapESvSYPeng640+vApUq7HEK
02hSBlgBLGo9zAith8yU+skfszvh0E8eFBWWIJ/G1gPQG4KDYtjEkl9fiy7tWTpzAH3LfT2F6Bx9
HzZUXmdhenrAtyC3Dlm3hj5A4pbXZU6GMh6DHMfz1QrBkxGpYO0MidPsl5fU4SI3BVgGkS+7pY3o
srMGgqQoC0fdxUCpnvPDX7LtapmGqhqi7r8OBLRKKSejN7g7xdzrY++TBtqGWATFYWCkxoBC/t78
QkNrPIdRQXz5ozsMdGqtUY8s0vLDib1yKXXQDlzshI/6MLxZhdJTW75Km1VOIa6gJ3DART5i3Dl9
rMGrPvSb6Nmm3hiRHBOf2J5Zh6StTeY7jrWuQAVnw40JHNNM3NAk4zF8nWEShyNGw4xvFtPGp86x
iNQXgB6uDp6Zzp0RKzDJBPWcyQaDzu2kU0fYL3ovdVPECSFswAza4/6qB4BDAtyauWScrWEYDy5W
zt4etC2bQZIAOoWjMBHs04wq7N8Jb7PWiScTTrad494QCTbcMwlQnzGYc64iNMJktOwDz4YLqKgT
kqsaCGGEFjl6+xUzuHw79+vJwRLWAmrj38Z/GbfOMT+IOMpGX8lgx4WTJoQUUTYXpB6ZTo0iaQTO
phuIGG+frUI8FOqcTCTUadY51pez2Es2eWQNBGefLRuDqsQD6IR/uKbvGRldjeVmQVRdF9qr4z/Z
BTR2wJwM9IkGdvUZQIFaNYwJqT5KFE/pe2tyJc4hM4016jTp2ZiT2qwrvBS6unyxxKdJZmc8KyXr
Nbvp0lfzRPvoDDfyYSbrgAZMcXO9v6iHNqNGstcyEfrZRqGH5amaIZLPk8Xch4a3LpFS76bKPpSb
0hg2IFZYAOwpVWESAZ57UMmMCLuncv8KNWBsGyTU3dNN1MxAfWrG+MK8XYbTGYkAL2r5YOXHelo0
PifwW3N9NdZ2mV1OGPM9+/YV5CW1+MChx44o+D+VO+xXhQHpA/ZaEDLP3HxIB3evS3uqKNm20xGo
cgMx7+UeACmiYANC4sZ5KSht/7stcVaX+AO5qhSw30jGnc7I30Dodx4qiBanbwJJXvWwfJCr6Ngh
6LWiHvcE349dRtkiZEFlq1jXxgdSTv0OLqgnvU95LqaepzMI+qh9AHNnOXaRwwpAnfKWYyhhs71D
bHHnncZunF2zF2di3EIE6KJmapNk3NpTi0o5Z8+aWlC3aUn+ke6QnO8gUPq51yMO+vVdD9c+RsCJ
0wFyvUFHQ1Jz0LVWDzopSPXuHxk8qdVsZ+PN4JXLeI7JYDlPsaMCfWVNOfqA5V7sGdl4CyiEeg60
iHQKOKUC78WgnnD0Fw==
`protect end_protected
