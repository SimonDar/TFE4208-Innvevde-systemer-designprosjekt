��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~?��^߫y!m��F���N�J(��5�{x�2��|#�Ήx9���V���(�R݅D��C���1��D����g�X�*���+�����C3J��"2���+x�$�(�A4*k�C:%��A(�9�R�;O 5�;j_��
�z�1z�@�����~���F�K��"}#�"O'�8^hi���k	Tx�UFI
���5��������qR�|p���q��� mQ�FSL��pK�?&T��"f��KʥGԦ6� �-��l�y��8�EN;��|\p�&�!�����RZj`7ZZ]H�l[�XU�������àx,�� ed���� ��S�݌>Q+�)��O�Q�aa.ߢB.�|��?�� {�UI��N�ޕ����۟�U��>��f�^wL�xLb�+[�ӊ��9J��|�  } ���`�d� �Fގ�ĩ�/�.�2�#���ͮ��n�����xck�(d$�Iz)1�~C&��w.e���w#�)�'�E`s=�Gñ��%f�;�)K�a��]AhҩL���잓��������cϵ/��:�5ԛ�l��ur�л�.	K4��#0>�%����,��[ ��G����4�\Vmd��=��5�_��"�$�����Aq|s�i������X�p�:�=v_�h]?{�����X����~>�[ ���<��d����Y$UnF���j��(u��6���f`;���		�@����mgf������>Li�0�m�:0+r�f��S^W��>�m�7 ���$U�z��$wXB�-%�D��r�3x8GrO���ek���x$�X6R\6��l��1�~(zޖ�V�?�����ˀ��ǻG�3����ua�Ac�|