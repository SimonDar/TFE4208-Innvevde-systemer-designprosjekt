��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j{����`�� "��g����^��&.���2e��,��Tme�hX�������x�
s�04�7h�ֳӮ?��K��	�!�n�:��YMv߁p4f�SND����3.�ے�l(���!�rS,#V��Ni�����g��ӎ���^��{�_/�0D� �i���vח�˘,�n��8{�|kR��W�r��AO߁.���Oܗ�x����~t+���W7][I`#HR�i�'�t��Q��<����U�XLD
I�-��$C���Ċ�V��b}��G��C�y2dle��r��f�%�%u����Ǟ"�y�Z��l,�(0t}�ciXxQ6��L�?UR�8���J���g��p<::fe����e#�U��7rq$)��J?����'�+ ��x����o�6vӀ.]ķK��tiI��'�\E��e��e���`{6�K�Nu畵Gk���[��[�B���V�uJ`J�r����<o~t�D=3s��Ojl�7�Hn�Z�Y�ڠ!L�)W�oJ��=Pi�Ɩ!����^��g�v�^�a�|槥�m�mv�aA���"�nɖS��k�t�����W@���[`R&�"���J_}��Q� �[h}��3� Ý��,R<��ЂĒm3��-�7��N���רTr6}��i�'3ۅ.Ň�����ڂ2֠�3�4���y�Z��C�=j�Uv��H]6qVtgZʊRĀ?��r��oi
�v��j�F�p.���o�f�^CBc�u���q�	[_`O�Z5[�x���o���ڨA��i�R�I��K�c��e��ܰOݪl�������T��L�;[��� )�����C���̀��}���j>:!�|���&N͔87%���sG��xiO���)Yc:筼Ep�r'��77<�Z��֩긥0TeTeȘ�s���]���?���ֻ�G2�����P@{���KH7���1�n	TWF���&�s����-o��Լ��n`ֆS\\������0��E ?�\�=4��g��^HY�A8<ĺwB��R)Ӱ�ov��zh�#�K�wW�|</���JpB���{ė��^e�uЦ�g+5���oatɺ
7��r���ߑ��
gw�tS_�}Ϛ#g�cz�u�
m�!V�O6����h��u��b�p� �G�#�\�{4B=�����d(;�8D1N���Ӣ7F8x �Gw誐Z=�C�'��r^}зX	Cr��hB�$9���z��ܠ�������:@�L�j�� ���Q�Z����/��8��t�iX$��Vk�­�4��H.��l����|[zk¤�S|[J}P;�
<����d���#%΀��P�Ed9�E{k�m��x[{Ç*����m�ٔӽqNj��Y\��]:���{2L��B5S
l���v8����9{���*:C�O���4Q���?��+Yg##������)[$0����	9����Y���� {s�������L�M��PHʔd4��$�A���ZweP;���^O����1"8#��'��U�t�`����eO�9��������o��ΣM�N�[L���K\8YtG>?��|܌#1�!�ʜ�V,RrX���:�-`�=4()�8�M|��&[�fY,�L_d\�+.��
j/q=�4�լ=�R�h�ү���Q';���A�ƈ��,�7o��;�/2�l>ep��7�)���G�}+��*�� h�py��gWPe�HD�D�J�����cα��C��uA��R�L�*��l����7\w��;w�B�HDN��-��醮m[��,2�1|z�/�)��j�TC�]ׇ>9�?Rl��l����b	�b�K6Wdu�b8N�2�>:�,�Ǹ�5l���hS��S�hyڑ�2�׍�j���4�*�Bۥd���x,��Œ�Ƒ��39>��9b6Na�H��J���(K�
�;K�"`�W�W�i�`�_3��:)m�;�Σd�����C�%�E(ۓ��� �+p.{@6���.6у9bCss�vrA�W!��
-���%x>�P\�����q�2��Zql���O�f�Q����D<֚ ��ǟ�pn��$U���5r*h,�>��l�%��2�($��}�Nv[E�}��k�<�Jƅ�2��`O㋊xl)��!KV(T�$``��n_o>�DK��e��c�:%ք��r������}��eX�w�&�A�>�9�~���֥�z��D��M��s���m1ʕ���-Ae�yc�5
��6���nz�h\�(�֋VKAK���J$�	%��)��r�Ǚe��{:��G"�0f V�,���8���q�k�]Z���;��ibU��^)�Y*����c~8� ��V�����*G��a-d,,<�gvA<o����n��	/�{޺ |���Q���.s�ח%���l�og�ʶ�b � �V�g�i�"*N�=��I���꿫f�`7��u[��]�^a3!���0p��y\9��IDG�/����^��l����a��n����@�m{�����a��`���2��?mkƏZ.2���ڗ�C|B�1�2���-�A%[P��;3`x�k�l��N��ۈ.����b������&����#�їakGD�ѷ��F�D�I�R-�����;l����|]ke�hh ��O��ßu�Q4����e�m�L�~��"��i��"5��(�8�W�6d������eAqPl��As��>���6��[W��# �e��Oڵb�-�bS�Cy��ÜX�cm�& I.���^��F��,6H�6z�)��q��ux�ߍ*?MJ�g��j�o�I�c��|�����'���N!���0����՟W�?��Wba4�uui����#�K*)��@���s��t,�tD��8�	���-�͸��?����'��=�˓�*'%=>"�s���;C���9Z�����xJ��R����Y��	�#O*0�J�&�	�DƧ���y�BǇ��r%7)����q�J˜��h'
^<��{@4��t�.T)ϋ�W��gR,�rլ��	���o��%$�$��L�Y�(�1F�/�T��ť�ށ���Z��ʃ��C���GTN���l+޸3	�1L^+�ML\Nտ����G2g{���%�{Cie������M����,H�Kv{<�	TcT��H�ʑ�\76��z�i���g��Z�;�%Ķ��Q;~C3�Xr��g��md}[W_+��4�&�c�����^��!hƁƶ�.p��\8Bztݫ۔c1��F�1��9�֤���h������Ε��94�6C�u��Đ�P�|����wĊ�/�/��h��/@�)�Y^��b�G�Gx�$�͈�����ԚN��x��%\�#]�!�Hy:��*&�����G6�i'���E� c��E��o�g�ֿ&'Ѿ���	����s�(�@�E@S��5�1�U8e��Dʩ�`��Ԍ��mz ��:XBn����w�B���De�����yrZ]�R���>.u1��;�͙��Vh8d@pzޔ�����j:��)_DI��H�8F�ߚ�����>jك��$����9&g3*cD�ЪY�D7SΕ[~����s�E�[>ѻ��$y8�<b�����������&C�b�Կ��;�Q`y?�V����?k�{��>�؋�(�Ċa�X��� �p`M.�����6��^�p9�@���MKW�1�Gx�IZ�
.W7�P6��1�K'�:%��2�I*2-�QD�^�i��cR��N�����@���o�Gk�G���6�D�o;p��r�sa5BY�bP��8����Sʙc֐1���S_ȊŚ�����6�Օ��p/ �3y��y2�R�v�Akȁ��?����N��d&����`���֗�Rf��n�]E_l��H���
�N,�V/8��pGo�vs�c׀�1�����J�����M֧��r򨃙��P�k��2[�������k~�俎_�岥,��
���e`<gy���4�mH��g3�SF�E�#�T)ʚ<([���,�(/�髧?$�]$̛4�|%�/�&K�8	k��d�5I+��2���E�L��F0�������y�K�|c'"F�HY�%v9McDA^C'��P���W�u�?m�0dL.��i:f�J�P�ΰ*ú������'Cnb-��S���䗈p����DN�-	Έʀ��ō8�7�{X�pe�6+`��}�H]0�:1S*&\t�������m��Ց�.(����E�~SS�YK�P;`��!&S�=g�����:�3 J��3�z��Vж�cs��*
ito#r�Y֜a�����.`��,�%���m66%��дT�h�4�G"�U,;�Zj���4�s������F�z9)�1v�E�o��%��K�����e��|�'}�_��[��7)��ڟiC^�ȘL_q9d��"w���^R�s[)�9���?����V����P���.����(ߏ"^kK��t��x;&�.�7 D���f7B�aG&���H��')'y�'��9��w��b�y�IQ<=�(׮��'L�T�$Wj�0�5�pt�HĖ�%�a��D�g-Gg>u�v8ɧ�s�^N��G�'� g��H�P
�l���(Ʀ>�n�X�����������S�T��и�rǘ�h���?J �\��	��R��}Y�%?��1�<�K	�X�1-)���R�}ج��<�{K����\�Ў�{S*�O�pb_��ު�nw�����?ש%]wE�KT�U
l���.ma����!@P�:�w��z�{#f�����X\����C�B�����b��wo�c�Oܳ�&g"��V�\��?�˵���=ѷ>^e̲/�p��L��+��TDJ/�HB%�1�]RHMZ��z-�&z��a��Q(u�DL1�������XZⷬ0�z/x� ܟ��������Q�}A|-��Ä�֟6���ӡ!R~��y���E��"�8����� �G�0*��� ����9����:����Pe}g���?I��"�o��1�g�r�u���_D1@��0`�d�
�U?,<���I���4P�t<�}�VC�R����`�a[�{�ྤL�uS��d�h�S�?6�~̪��JA1>�����5��e���
�	^`��1'&F��z6Z$�xc��*�;)�e?^K�M�u���މ?�g��y��{��K����U.x�ó�	��	��"��1"l���������Oc�f-^�,�	�ܾ��e~M���B�J����xm��m≈L�m�����k��99�b��U �C�l���l�bv��c�LP��������TZ=}����D�@��ܧ��V��!+�t�{�e~6҅�"� V�qv��`�i�c.L�ax�4�+lg-H�r����6��(`�0E1B�n����o7�)aZ�3R�E��C���0y.+8�ܓ|=;�x��]���m��H�k�D�-�
�6a��j��� ���UR�޵LR�ߧ6��/������A����2�"��G�gAL����djm�Ld�_%&���d�g���R��A.(ъ!�9ľ�&6��=�T���h��r�x>A�t*z�R����&��S�o�Ȣߦ������e�Gr@��X�4����X5��9��y>���t����L"����i©�� �l:NnwHLW�i&L���]�ͪ\�Iٟ��!��^��K�o���"ǫEvLw~�&��Q�F�Z������i�;���{w吝�a?�0r���J斐	�쁁��X7�ק"KC��e��q���r[",���3�(���**2vhP��B��R�Mar��N���CJ���-�Uo3KDsN"K�������E�M�`�~��q��s��[a�\�>�M|�X\�x�w�[,i�|Y �^���0��L���K5���������.ڜgYn�y+-}� дu��MC�ч���	��u��It&JhӾ��0�|��j�� 2��j�k5��m���t���?(�O��q��� @��� �������P
����-,��&���b̀��X�M�2�Y���&�������v����r�8��N�H�D����޳ ڒ�R�@��?.���w�"�@��7���1�-Ma��&��ݵ�b�� P�9�Rxaݓ�'�Qgؽ?��|�X��~|҃�6��{1����a����c^ߢ�_��>�ު{�#O�t�C������/�p�βFȥ }��ߗ���5���ԏ��q����_q
,4���`u�bK�S��OsL������6h�ħ��f�����Έ!x�i��{�m \�K(1{���?�V�r�VTqyE"�%�j��w$�x���p�M#?�W�3�ʸ�z��L�6L#|�-�>���a�B��Kݑ~��oA!�������J����|٭!>��Sg�p�?N�_i��o�t���y���n�Iu:Bs�CXq�0%��� ��DM��rچ���?StK���xd�!�zy���l���,� /�u�ʄ��f��k����'��KC������,H�x ���+z��qpX|L�p)��K��fFi�P|P�>}��31�����V���=o��m ���='���)�8k��;�"c���'�SS`�"��I�`Ӂ��Q�'iߴiN!5/�[X�l�0A�޺�nL&AP��g0T]5{���-GL_�����`��א��5va�=V�襈ʅ1L&�e��ywW���%��g��;�$�В�	�)J���Uc�2e��-Of-�`LYŻ�$8f�#o�6&�V�o���­�7W���0�xf���n�:uR#�L�������d&܋�4s��}�;S^\�X�����.]O����F`�v�گ=%O��+��yT�L�/����~&�Q��z0�_�g�3���t�L�?X��礧59I����{�M6G�G�@�ӓ'��TF�b��^��0�ٌ÷m�!Y� ����U�X�c�A.����tN|�_؝�V,8Y��7�M��:��b�����P^~��),�.�F�)��]H#��3������]by��C|K�8��|�pƚ��5�\��%K���O+��r��W"�:�MѤ�]F/���� ᇲ�6�ʙ��������P����-|�e~I%���C.	6,��8ǃy��O��z���$��ΟQ�t>��X��{T|���;�m�iR��t��}r$f�=<��cP.Z���⿊pĔ�8�$RZM�t�fu�����b�+z:_\�z���,��˲��e�P&�\:&s�����uf�]R$��<"1�Y�,�����s�� ���&;��H|h��nm����RǮY3���Y
��J�����D�%�5��R?����od��Z%���4�9��m��6�k�+bF�~�lA��*ƙ��a5w`mjz���|JRl�[�-�k���G�Sd�c��ݎW�}#�Ϥ�ۤ?�A�#o@�7��΄�/�g[�R�P�x�u`�Q�~��2��#�䗔��㬶�\����s8���[^5U�W�r��/��<�H@;'���NG�I� ��'�K��AlI�)vU:^ͩj�[l|�?1{ȏ�S�$.�)�ϸ��!��L�]��/�9�+��'��IC�m�q�%+�h��Y�?�� ��@�'d�<��V��*>�Ͷ[��ߤ�X��FJ��vW�A0�nN���|�.����[=��N�ʀ���d��_<0���4�l@�^e��*md��`}��1wqs��U�W����+}�ß�잚&�ܾ&a�KM�w�j�c�A�V"!3HƢ��{6L]ўH��b��'ێ����%Gռ1pY`����`y짳f�+K'�Df���.p�*��:�-nPRr���|L��+p�pWO}�D�`����VV;��S�݄�H� 3�s����%����(�܅-����'�������?��D���)�^�-�a�VՑ3uE��]�	�o��<pq&�� 0�C[U{��o�p�)�t����2Z�[���Z�t�I�I1���E�	ޓg�Cq,�E�XX}�α��z��r�qE��PN��F�t��ݸXU�F�P�����6L��l� �k���N��� �4��I����+���0%�$�)R�HK����#$e���M��wE���	~��+�_��[3�߄Q��0���Q�g�f��%Q�B�<h�D��A���r��S�+�a�L��H�@c\_1�.�A��7����V��mj&lq	��]��bB�@�5��/��瞵�Z-�Z�� �*�,��h~Bs�����`�ǅ+{�@ G䤬t���,�=�X��_�{"�o����z��/�*>�F���!MJ��خ�|��R�?B���ܻjˠ�2Q
@�t��Z�