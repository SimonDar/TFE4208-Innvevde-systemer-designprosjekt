��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_�>/��zTg��P��Y�@��+����t����m"�Q�e���VW=I��K�']��GBI��|vz�ٸh��?8�2փ�%+.Ht���Ĝ婒e�])�5�Z��yRUn�M�����Y�?�8�>�R��2%��y�� �%����*2l�o$'6r�A[�q� ���1u�Fe���r����.�d��@Lkc���f/ϳ���ZL�|(��o����:���D������޷3�fiq�����IM�uw��xC[�gK5�ѧ�/t݋�os��f����ݧ��^�c�<;#���J�o�
ͦ��!���ˇQ��\��A�Fo�؜:��f�)R�7B�E�U�Q��T*3o���1�l(�bs��X��?�ڍ2��,u�c�͹��܈ۤ~��:�EP�h<C���f�̧�ܻ��� �cAj��k�Q�ݢ�O���F1�RAݵ���7{,��[q�>��d����j��������X� ��V9��g�aT)�T%�x�)��1V�ET�����vw%uX �~"NS��=�IT����h;��<�)��cRz�oQ���m)-���-8��߲h�l�A�r6�H�B��/L�*�a 4h+�:S�"K�x7�O�Գ��_��Y��5&j���2����2ڿ��t4�M+����<.�-Iw�˞`�J�^;D����5��)WT��|ɼ��A�u򚡔�E��@��h�R�	A��*_�O;U5�n$č�xE�x��&���ʕ��4��i�k���_�s�k3jQ��ps���Z�;�N`d�=~�7R��F�$��ѵ�՛쀐m�u�� Z�a�	�ٌ��'�j��[����,��EW��q�dQ���=Mج=�+&�c��:����~Lu�)�v�"C�� �	���g�A���ؑ������⊃Y���2(�b����7�<)�}~'V�UȮN�|�q嫾e:A)LN�֕��Nmɷu����US�aC�;��|
y�ipx@%�vq�-,v�fXekM�b=���l�SOD��.
bs@��w_K@D�D�+����nȂ\C۞�n*\�X���:����JH�[�_���CĮ�J�s�J8�>��g�T��P�)�����p�N<��5Y����}n�W�9$��h��o����佇��'&���g���AU�/R��q�ԍ�]���ɇ����B��;neԟp�OXձ���Ye)ߠ������RV"�U���]�ȮɊ~�v4P)�]�%���0J�+�1]n�ɔ&�m44��{w���yYEϐ��L��8��H������>7��m+�����c�*���B�ˍ]gdf�(8*��K���̩Q�ta�$����Zx�{�¥y�q�ZH"~�0^_()b#������I�l(=��5��Q�P)�~�۟+�L��֟O��3yʦ��!l��d4t@�j�Mc�H�o>ǧ�/b��.�\X^� �&"�G�vnm7�?OQ�%-F�t�k�k�-��� ��+�M�l\��8���D=ۘ,d;mkƗv�U�����Cc�s�7��'/8vp,���`"LKd��q��Y��N�r�g��k*Q�ժ�Ֆ\��ǜ�Oj�R�8:�t/M.*�XS�h��A��i4������1�oݨ�~	�빘'��0�?C��=K� �,�ܚ�Ϩ<U����C�y����v^�nCV��eה-�A�'�4�?�}���IF%�j�TkUr+|c�-ÍQ�a�@s�ӑf��}s�]G�4\�=�\.�5�6s��� ow�,�1�rcX��(�z������>n�	���=���ͽ뾦��K=��C�J�W����9#H��"��
|{���trM�Ħ"�j8��bl��L�Vk���!9��]�i��g��>��o2:2���9��g�<A2����hd�]�zq+���Q���u�xr��.�c�]��Ri?<	6ݐhP)ďd܊�
���[n��7������]���V�O>:��3�*�'j�0h&y�!��M�N=�z+�����T����?_���\?K��(x6G�ȫ�7(*��{���\D�~?3VDދCϑ�c�(ϼ�t5)�LC\_�b.�u�K� 7,��Œ�v��j�}E���t����g;��k�1��2�5G�^>_ޚC�X���~~+&K����M�(��H��mIqQ�wVJ��=�+��4�k�^�G�zd�Db% s����[d��0��<���I^�]��p�W3Ma�k�S�}�Ԕ:S�	M�^�Ƶ��^�ob��	�TM�͔� 6�?�H���޲ձCQ�졻�4�'W$z���/{�/�K3P����V�ܚ�������O�u_����+�A�B��Tk?'I2� ���Sd7#z�)�T�/hy�
�eXr=�6t��T�O��zQ���6&�����M�$P�ldJ:=���?�����~u�e�vE�<���r������Ҧ�X���o����|$1P��	��GA���A�Z��`�m���"��W�8[�M�8t��>�����c�m�R�����7qL����~�A�/D�X���h�&����v��jo^�J�R�B��0{L����� qOD�p�<����,��vu�7�Ѷ|n��:b���'6�	t����q��w��4�/���Q���ǅD�Xڪ�׈�{����<)�k��NF��X���xۮ���扝v"̕��}���bp��M�:�4�/0�'���ۑ��̟�ͺ���9��3�	N{I���L�'m��p KM��i����`�:���p�}ҳ;��`�-g�e1)�3�.�Z{&� �hǪ�u���;�.���;-�/s�������K\��{"gKv�px'���%��/ d��`(-��	��J�9�I�#� �%¡�&�ßt5���6�?�/t��Q�*�W�=��~�G��U��\z7 7B]��\���3���u��r�-����e, ���L���?����ɣ_�IB�.0}Zm���o�A�ʻ��C�ސ�%[��:N�'���Q�-�S8~A`��Y��`����=�� ڍ~���5��޲�Z|n_�%��3A�����ZӋ�=��,��D��p����[����c+b
�,̿�h�K&�@s���K����ҷ��1H���ӽ
�2�D ?Ԃ�1E��r�>B[�}|\�E�W�0����
R���yO�R���Z�aT�@�tD�cF���/7
�&��U|	W�5�fg-�o�4y�d(��K�LM�ZZ�*��B��_�N�o�Y���9C���_��7=M�d��Z�]8�(�^�
�R>��W�2��|r]?���-;��0�#�o�М/�����N��,\1V��Y���<!��j��v������qO�S��L�{�ܱ�I
K#LTe��Dʲ����IzՏ|���&8|Z:6F/Z"��l�mv�7�P���V�˛�&"�yG���/`��9��qM�� ��g��������%yUX�d��a�Z�����v��z�D������&�*�Y(#�x?2�B&�����HL�TU�-kOM���i�Aτy���	�g� �ѩ�BSh"B^�0���$��W�)��	0b��ߋK�ؾ͝���7|�p�(9t���{?Q�2��J^�`Gv�U��#I3����8�~��%o?�o����x;��U�3)���6R"܃Ӑ�_��4:
}�z(����١�zI���+}b:�x�cۓ]�y�,f�T���#gT�I�x(��@� S�D��,���foo"�h��&��#�e>�{cN��G�� ����m�K����`�QbwV|�����}.q���7�eU"L�k���ƎTw�.�9a\o�ۣn!Բ�$~��{^_��ةQ�����E��&|X0��g%��-�FZ�x� �����W'h�Е����6�� p'��Qئ�E��L�4q�}6�a�1R�7	0Z}j�����c��'׎��ЄJ'���mpWy�$(����(�;މ�P�zcP��V�ad����{�P�'1��ñr�4d���8V����"xz��.ncBc,�M�_�CK̜��=��w5�/P�wۉUIM-�R�9���)�����W�R��_�2�W�*�gO|����0I�P��Mɢm�g�B鼴��]�e�ȮC.�L� �6�aM ˇSnȖw�OƂ��Tp�%�����{C���DI� �S 5��I��Uo
|=��^
�͵�P߷�.��Zn㤕�aZ�rǆ��vEDG�3>�!˿K;���׆��lZ����?���,������Zx�z�t�)b�g!B�/��D����=O����;0 �i��gM���Ԡ�ă'q�	y��kwo�W�<�g�B@em����_$���8�o��9��Xl�������rz&�>=V�AIp^N���� ��U���tdZҊ9��5r�e1�ب��E�l9����4�[.r�#Y��"!��%���P	���m�w1^�/��(��D^L]0��)�p��Pa�Z�D\�Z�0;��ׯ��'��c�@kZ�]�τ��3���t����\��_舯-�1���!&J�|��ר��u�z��Es bD�"�Co\}p�5ֳ�YSZi�|XHC�U�me�E�u��_��V�C,pk�g|��̫Z�T��:�1;���#������Ɂ���=v�~�<�d���{de8T�\µ;LeIu�b俓{�g�z�B;G���1��g̥N��h0��1��O���VNW�sIᖞ�y��pC�
@�Y>��	JS��P�%���3�S4�T|ll"��X��.&��Q
#s���/���@+�k� �_���4������C�S7a:����>u�O���?X�6J��mmk*k�a!���&���2��C\�R7�$ ������(���$��|���ߟj��2do��l�s�L�(ȏ������䣉��6�$.�|T�vq��y1���G����x��,
����Cun�r:�K%갳M���k�̮'+�|�tmAQ�V���P�j�D<4���*���3@�)�xDI��u��:�#�i�T���D�v5��Ij�j��~~�Y?jqFm�/�?*@h������hҒY��<�"L�s���u�S��|��2�	�b2��Vm
̮�'*��"ס`��u1��q���BB�S��^-���W����7�����Y\y��8<0�U�3�k�$�S�Gd���H�0|��Ӫ��O�r��'�w>�'�3y[��S�v=��v����!�ƌ"&�1ok�p9Ό����ة���\)[���(���2�V�x<:HWX���@��3ަN��<�TS�2$SK��Ryi�2���,��6݋=���6� �պֻ|�W/_9N�W�;��?��h(��y��oHa)jTC,X�[��'�!½4$��g����?%�A�P_��
������$AcR�!=��}z
X�"	��my�e$%F��sU w�Yγ�z@h��E %a�,�Ƅ,��Ć"m�j=�Ys�%�I��ه�i5�\�Gr�L��=��)�&���<����K햰���
�G3U2��E��;���X2�.뚢k�7�g�8����t,8��?���DjS��6׎xc�� �ni	U��m�U�#�|�3���Q����쒁
�&<ȋ_0�$j�ni��u��A�T �s�凹xE��������8�:��~&�CԮ��mt�N�A�N�U,B_����î�Ʒ%b�+����Qq?7��&��AM�u�{�c��I።�Ҷܪ��oF^L�F3����T�aρ�׽��������7f����_�����Z5�UҶ�څ�����?�ڋ{�&J*5�3x�thz�(c!W�f����V(X��'!�����U1�~�Κ���`��=d6-�n7v/��6��!�Z�U/y���M ��1cն�0��g.��S͜���&��$�)u�������U�q���ZP$�N��H�~=P�d�v��D&�C%���@�5����8Az��1��W�#�;�i�$�����Ri�!�`�4�f0����0|��h�PH���ܢ�~4,���SS���M䳓)N�v�&;
Q�CgV(���g�v�>l�x��)ct{���G©� %*� ,�"� ��K�����|�Q����JrNp�M�t����Q�Y6�d�G��?�#􊮩C�xM��Q"�� ʑ"����<���Jw�k�]��*u}���u>m�CL��2�B-���ҙ�¬�� -���K��Q���B��e�h;e^ǂ��-L��XM��~��:�i3��s7��Lf: ����$\[�rh�d��^QɐTj#I)�����L �a lA�,� �&!� ~=��[a�<7)7 Y�o�\�?s�}#���eݛ��P�&���}=ԧ_���)ײ�Q���O�C�� ���d��syu�삸��R��g��}G��0����ObҬ.��A�a* ��y�W`QY�,)jw�����3�O�Bjq�`~ \Q�:�Ȃ+'^vW�ҘƁ�SR�~aNV�16�yp�H��޲�=r=E�4p5��;$���Ly�ᆢ��ve�fXJ�2x�X�P4=w�YXj"$fL���,#B�da��]�x<�>�%}r�����#�!���Z:��Te|�y��t|�0D�����eF��^I���։E�����j"�f7b��L��J�P��kL"�����澯4�>N"��yX3H�$��=���^��ٸ㏬gߠ�����@�T�
�]=Ӥ �E�;V<�b4����P<'C�A�c;	5)���E��NIVϗ>#�������CM