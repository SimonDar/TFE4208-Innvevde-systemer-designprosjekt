��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�I��9���<	gG�����0 �)���*�:O{85�L�M`t���7Z^�:>i͡凿EƧ���ڨ����O�&�0j�u���ge��� �����������W}��P��R�<g�����w�O����]C'�N��B`��ρ('���Kju 
�	��Ҹ����7�#>
�����J����C��6�����`�Q�\��xH�xyxZm鈠>%�M�|>�L��
��6jN�b|Ck?�
�ɀ��[�"&��q�X<���h<8�$�q�o���,�'��cf�P�,s�����-Bǩt}�y{X~7�Ȑr���`��r�-G�/���S�wy�Ы��xՀX��h����R��W����WZ�ӣ��fUU�*��2ü�;z-�X�ub� �IO��$|y}�O=Bwvv�����5D�ow�a�w�v>υ�8$��M�����O`�l��x��Eڰǟ�62�z׻�Ma4s�8�ut���l��ؾ��OJ�
�GMɴn�4��]~�U��C���<@�e�G��]��T�5�bLp)�j]Deu�����#
��N�:��%$�~M���G!��<��˵B%)��"��6�����굒���l�,���/�.-�(\{�T���F��8 %?�:"XBb4E݆z��\��
{	��.���}�e����R{�� я���AM8�O]&T伶��f{��Amf3ji��4��DG�b����ili������ ��l��TEK����?xkM�A��E[�4g��{�F��8,Q,΃�5p�A�,p���TH\ױli����v��L��럍��4��8�?{�b% n��P�#8�m��$cj��jc�Fp���P�w8l��Z1�"3��~{��)V�ӰVIs��A�D���+)D��+I=�/;�4{���4{���D	���k�m�ϝR�������?*o'����v��I�-ݓ�QA�-�J��2����\r����l�Ly��w���M�!���y�xrY(�_L������ԹhP��-��&�*{s��%�F+fjv��W�ڈTC^.pהh,T�.[e~����,\����ݵ�70����jSn�H�e��Pa���V�d6�������!�{ Py��\s)��(���@0�X����=�p/�|��D�����t��RMC�&�w��^�D��$FNT�q�,�q�#��9�f��dA���\;j+��07Z��|3�
��:v���^x.L�d)B`�;YKy{���y���a��lס+���fa��Bw�5u'߿-Gf�Q��{I*�$Z�:�F#�����$�i��^������Y��|q@�J/�-��v�<�p�Ƹ�t�O++`@{|�����b���i����p�_��-�o��NKO���"j�|���z��<M/��,�:�-S �ϣ��9���A�T�W�i�wXXSӦ��Ld�״�4Y��U{к�V�4��%lBev!��$j��U{|�����mNcQU9�ٝO��C-Z�GX ��y��$\�G`p����V�����Ɨ6�pP��J_{j��|�I?�-Z��ؗ ����(��[-��;^{�>Y�p��#��j��f��'�U�����Y��F�CG��(���OX!��2��j�d��ض�F�;�2�wu�&g0sD<��ڢ��Z��*�?�R�lꊭ��x���/H�"�w���I����K�E�m��N�c 2��XU��/bG�\57_Md�l�o�vP���_]���3~q<��il�5��	�J�+���6B�]�d����_����f�R�6��������?��*�˵a�ni,I{ ��/��e	�ENUOik�.�]a~�X��硲t%/�V��E��F��7D�������x��B��݀%Y"�&؅��s��.�D)~ٗ�������r��/p
���ޑyl��ԫA����W�fz?�+�0\���N�5F�r~�h�V��Nb�i��Z�����P�SW\���Sq��t[��(ש��̝��}�S� �F���j(=M�c:�+��p��D0��a�qܑ\�N�*Nv>#c��HH�ٽ��M�m��0,G�[�M@~����5���^���V�[D\2�q�\LF}R�n�n�=�PZ��g{@��B��~�=����iP��{-�+�]���wH5�?���K���=+elC�0���H��g�=�3a�S��`F������B�_�2�����]�_��U��&�c��/7������A_�|�+/~r�L^�ѡo;�{y�ḂfG�4D�n�f"̯c)֋J=O����õZ,���i��¨m\`@q6+�	�+>��PE�G�1�ٺ�
q���7�oî������mR��i�g�iǌ1	��<�߁R8Ϋ������jd%V>}�nk�B��St+\� Ɛ��K�?�������	��%�*��L6�Uw�,���{�L��(gCQ.�T᪁W��P0pMQ�Xk����	^�A� ��}V\R��;Q[�"4��J�����ݘXj(�����_��NlճVk�K������> =�ʼ�PL�܎�AI�>�l��&-�~��Q�z�.�q̎!a���{�:_������6�̏�5LD$�؝�Br�`kh@���'/��dy�F��g7~�oO\)�L�W��ޞ)i�\�y���Ky����?	�ʯ��\c�doW����J�D}��X���.�ad&Ik�*��M�9r	��l�����d�1���%�v��lϵ-^"l��ޅa0p1˚�g ��j��;R$��\SA��|M�����IS��`�S1n$t-ή� u�#�ϰ�����[����)f��X���̊�F�ok]� ��=겴�	��V�)�m�o���3ǟ�Z] �C���VϢ�i`� o��2���FҒe�����T�F�C�yq���<�^|�L;	Z8�.���Zʯ�F��	�K�9l���Di-�g��u|ǋ�F�o��r�\&���.h��A(&W��J�4jZ�=�J Q	��v�Y�B@t�� 2{UqV�z���u��4V�( ��M�������ٺ�fm�ъ+�.��^H	NR�ex&/�}����Y�ũ`�����t����Z���LDi���R�r��IU9-�ߓ;���
#ad4D�(Ҧ�B�^��1�]��0r�&�J���3k�l[S����ǚab -},ޔ/�:1?$(�E�`�ɶҶ�������-�W��ܓ\���nww(Ԝ���*�6<}oUU)P]�`g/[��}&b�-R����\�&m,�"%PR��e/@�%���C�ب�_��s/o