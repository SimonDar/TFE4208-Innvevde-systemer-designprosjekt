-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
imJKX+jJzDwg6+LiW0ARMkLbPMiC+FjpK/cdwqVWH+nU2efBS163Ap0vUm+8EJU5jilSjUhx8kN3
o/cztAySZXUmRg13RejvZmXXYN5kkoLaZc6Yv2mkMtYyf4OgtEU8JEW40r5OGtRDbrswoRsSMQ/5
Nu/nTvRgYFSuJ9vkA6dQgN9iadNmQCEHEOoyoR5u9VkGvtdvCD09sF5CUDg+HxtU5+akJXlaRNq3
Wx6cH5tzzjubIMYEFSZ/TU0wdPTsGwvlyNUG+10E1yzje9hl4Lagk9el9mUOU0zNU+0vldwWF5yD
D7nDd9t1LdLrDgHZBNg39RNttNWRjNnCOFbxAA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
5Xg9uB2cE7Gy2/nN8On6b1h7MQgOqe2JIpNTsYg8Nq0G1sqNbI3wnO+dmjIs1SmLi+bgF9z2yow7
bXGXF52WqZfZmcrAMGRyCnFpEyKio/HF/FDKpp4RPdNMjTNVK8vKq0g12KAFoAt/B7SBWjdU80UK
yBWxTQ20UkmRbxgzG24im7eZPHY61jTzYFJBN0lVTBHv2sBAivIy1XarHT5KvhTjn4N+/zBwvY5d
gBxjiHpSkR5jP39SjVOqEqWh+H+Y0yCeCD1LqK38j1mON/B7o65lsiCu+bes1aygICGFLuTlb8QS
ag2uIZkbY4AqFG2I5ETRHYmTCcoSCgo5ZjanGONXUWC01kfiMo2/Dv5BQGmJ79WroQ1crDqCFQxH
mOh3Y4KDD0/Hucdv0z+QuaO3NwZOz6PGvhv1ipV6hLd3ypZuxPR+lYGS5Za9uS19hsCUVKXmzS89
6Mb65M8Eoj0y4CXmvYAKc3Qqp6yGsDH/ofSIoyilMFx9Zz3vRANyld3eH5lAaCwl2I+GF+V9ofAM
guevpUfe75K1WIgW/2Rs6LCQbhvG1C7OwwBTZulzwu91qIA6lu5dBEkpFFgJSrz1dLfPeMgqs/ui
4VQ2EJXBGbguczbeyjxxS5QjRVnbAoeELiR+CVjjW+jM0CMo6Tt+dVlxBO/6w1EZWPfrwg1xyLfq
QxS4ms4PELTtsbq1arX5Z2P0dTvQ4uuYiBPMgKTmO2iQBgO3b+e+wD9sjo8mgQxytZCAIhXi/iSz
RHQqqzwOywgV0mIrJrcTyIsZj7ePJnYcb8C2AqFklW4qq2LVFpbUpCd1naEQwRFh/xWIviSOkt+W
ZK2odaujtt2ARHYofproiLDheHRkhS3xGaetBlrAOtp8AZM91dur3apDjzYPQGU3IUvC1K5WSFzL
7+eIAhA2B0FhVNJEMqzwsu0vDhB8g+db2nac8lJ9ha6yQjSbahGgni1vOoOqHoGIqTUrs+NLoGgF
5tULPRAuPOIQEFigunrge9GO2rVlvldCwaYkMcGlEuEgzKtNG27uFPyVHSMFeiWsMh/+nCoyIvdn
EMv2OiAJEPHbjf4aTpxt1ZyLlsDFf2IyR1bym+IMoC/H6hFdp+ymV1yDkPoZ1I2GqNujhgHPqUsm
9jqfDLuv3+KbGvbK4IHswX5ciUlci3usnri2iFfKzPS1f5lYOpp+OwpEHLUixtRcAxo3UdmAdOJi
h/Be3e7K7QplldZdCiWEswa07BGOECool2WeNo6ZaZEmCge/r/Ngv1LOC6O280cAJ3EyBoac4adX
dZdWlvLhpNnoDqsNiEUTX02v+Y5LTrsdCG5ndiTvxWyyeEO1XIZE5UVjYhwKKqFRLmzvWUn+XUBn
deJmUoEko44XnENtudvXtHMn9SqbLWiGOVJqyVvLKuuMw+6J8UBlVRUl0Y01i4rWWg0983ijY+Ln
3e3pyYwMeTnf0af3HDLbjAuWh8Tl0VbHMPN8is+eBGslo3t1hIYKKGBs+LwjrCTrnmgYQx9Fublc
TqY2Vk3RjJvVien4404IphpPUivANIp7yST4ZaSCFtu5U46+ttjEafK75zTleOs5BL+jKudMZUr5
cBRji/4EBAJNTGK05u3XPjuLj4Oan3X3YIHQmMkOWrqsmd6facXAG5lhmOMs95omQulF23v5mMfH
mEayZrKik5RWCtsObaKloDNS3DBgUr3scyeQ7Bgf55YtlSdRiaGjf+uId1AoXuht4gpa7q+4aw48
zyRpO2Kiw/34thP1DUKKjZg0muAYefPzcIJCDWaTDeYLYp2q0lae8D6U/CdIdgATzptSK3asaJf4
uhlPIurEG5QvNWW30p2fjXQ3aOW1rYkQYbzpyzMdGMUg7l18MhT7ZakYZPNdwyuGs7e4gHIxMljw
fCtCTYJkeg4GUDUzATZzlZA9yeLbybXrwvJ3Q/ACg5ABuOmJiZox/+/I+ed6Z2ZAH8A2cvBSk8Dn
hfsql0SsmeVCDcvXg1zDxMFctYaAIZGyKvWK8BT+NBAgSs3rxJ7wRkag3N0gx93YXYMk6d3OloLx
zPQxFPv3WofmWHjws5WbTbWCDZ0XM8KtEr97tH9X3+lJtt4SuO8PO+16T0mcrTG4R72k05mp0iAe
jkGWLYHzR2uz6KbOZp98kQEky8BOlKaCkHxFv1Sp+oWJeox42EQ9YmvyQcfMqcFmWXXphsfdwFio
+jPl7UhhxsE6j3H0ubYpdFbR3mbdvCu8xH6jkC9DshE/36pnPFBHjnZkcBxpHvFKLlXNhkYeYChA
gIHE3m3Cs8QTLKb3y5dfM8jtE08xOjR7hToGytwDfzl2NGvKcUHEGkiQUJUfMzz3i9srbFC3q2z8
lZRZq1YoHEdsuybyExXqLhy2YN7jyrhwMcEvabKXLZjDZQVxDgn7S3IbAM0SuZ/vez5c0VbOrB4w
EenKdXBkLGrMQgZl2VXcwvDetxa7gKRS5h6Sz4vQ/I4WM6s0h6awGiG0WortQj+UeEdWqCDlzxG3
Qp1SEgbNTkgoHYsKmUXUTXjsRKV3cNAWmJL3YV2CRCPxS6/teoV6G4wtwWQWs9IlJ2+PUUlUIXUY
xrJFkoO+8C4Zxu6s7Gp9WWbGv6ZKMJzD0NRTKponiFzA0O5TPx+HrmBbINB3+ucQT83ImN0x0Np8
fWJoCVm3OpnmipiV714Q2aU6PO8+nJet9JPmj/s8gZPF4RK+moe7GbQ1HcW9E+l/1/I8F8he6R4P
e98wZnBQ6y4b8VTGMSksm5vQISF0Lce28xRVCiW94BexEUZU1XLr7TZPz/DcWjI89y2jI0ZF2quB
GeZXIryFp+nn6fph28WYru6gch/+7ch1ICkibduitVfX6HgYpNAHLRZsWOkVhJzkygl1XtsZuIGD
daJiwdup/q1ZDB1V2Q0cclTacFboPbc/HV8/0Mt/zJSjPYUY6lVw9axvgDaPi2HPCjj0NV7yXYZ+
8ZxfrIQZFPiq/TvguKUk9414GzMjFl9fBtlaymnOYhLsWHTbaJWRCvcKeVnnoV0KV4n2K2eDdMLZ
GBYLXqU/f3EVVU8BNohkkZJiKYBi9bt2ImEA/DM+2awp2w9U4IRz0v4aF3wDcqqG3cIg9+ECys9r
jKIST+hc87cg+yPWmv4085fjEKlx3Xd2cXHH9a1rqLYnqaqhf/ntDWQP/3hvezZAB5y9QUC+6/PC
uTqbeFQGj09Y6LfqxPofOh5m/mcugD5AQubJm3NKphzQwfABYXR/+7IzEYK94XIGJBqRG2stmPpp
j52cRE0HgWB6aVV7M6Ia2NCU44C7v2zaw6HBkZqgZ8DiJ0jIedV8gOp4BYu3M3+qCqu+j2Lwk9U1
LJEweWss1fWNgORDpbzHtXRJ3a4jEJgE6AGGYGX6dew5h1AjtKg42AJ4ATr7c5Q11/0sj8aa5BBi
LDBBbUiTLfarNvrT6w6ssyiqn5MUTPgHnwO9OJeE2vMNWIxxk8pluAJpMPQVyJ1NlWidHQIg2E4e
Abhbs0Ck6ZbwXl+bkc1IwXbPHu1pz6GehYRHRPhkbevwRguZPZCIQl2+5Rz1OBaHDzBGtI5F+3rK
p6Fx7HNWcwSTrWJdqcSyS1/q42rpmvT9PkOpvJcg1p5mXL5C+1mUz+Hdasn+rSbfYWmJPCNJ4kt+
T+mTNvsYNqPtsP58LlgbirT97zGW90YX2ZbrDiIJAytjgFCM7bIDm5fhBWf/am7f4Qpo4HfZgBJU
tRx3urTeD3PWYioBXPsf/a4s1ASD9OlirbagTeI5i423HZ5IXcI1pYeX8dgiPI1Q03qzZ+jHpaX3
vrb1UGKJHgu0knCsyJQAy29EsprUeZgdIOZT5EC0SQFW/saTU+l1IOwuTu0OnLTdKY/pK7aD21jR
Dtw2pU1V+yCg9eryv6eb4pBUlEjDKhN4+9xq0IWdZWaq/eHbb9jf66GdISS6Sdbajwydh+r+2eX8
LEm5ZCJ7vG6LBXxs9QU1cAjcUZT5mwvPJ5KRmoXdzwhF94XBMUEiSOWwX1X4RAiLNZwJ6dnZ6t2Z
q39cxnZN7PubdaIbbJUwyXJ3G5MSo5lfY+JoVSw5McBHW2cIrMkz1qpx9t9jYC9jLafrpZApfGTw
OuVHf/DP6u27YfHhi9ZX+FtBK7ms2XHuPDubfGTTjc6ah4QGyEqloCxwGHroH4pS134DU7UTsDjt
JUQPioCyd2zpb4dg3oxk77sbiFABU6JQIGjM7d/hcTIub9lOAkN6yX6/aCBwXgOm7WcrdoOBaUdQ
d58I108qKOmQilAP2BbmCz8TzYVvv1Q6kkFRSWuIQR4sBiJP1EXS/lWWANXmSobyPlE/eLEjZJi6
aNIjMH9wMFoYr563vbut04VBimwd7cYoI97JTD0UjteFxOZJDxY76oXMBQWpCnTrVwrA70E2TX1d
Xy1mg6weyd5U37K91tiv8zDjFWFaSz5TjyeayYBhMUePwF5BkKz5mdYkugN9SrO1i1e8RmeWds/n
3+VLs01IMzJ8Cb5lgzPRT4UUlqgIshc+0Lu0lVOedm5PalRF037WmVozpY67qE0kpQubJIGzLb1M
2GNCrnQZQ8axsH+89lZcfyA/ImfUxLORWtpjkpQeYRDTC5YWqiMTuoh+b7zYieN4j6sJ6AGpw63U
wuEtnAktLMGVT/6N9tSDcGzYWdxxFcwSmO9pTr4Cf3dqiqTvVvIze6GHT5VfINor5pldva1Bvs0E
lCLFK7CIa0tcgiuFSwmJX8D8KhN8EPi+gnhtljxkAl6Mdy4G6+zZkvnls9+BqD30D6EnEvgLpiet
RtZYxMvUjbAWfjAqOTMcQbNbW6AhR6mkYAtJGRzx5Pt1TL/pKOpk1JrwGzm2nwgoDhQxJ8B5nj+Q
DNXyTi8y3G2Odu49DN+NTlHVGvYU7NaZhfOAWh5TaHMhdGqU51iklVSO9SwCOsQhR7x/1z0BHtHr
ojBveDvsd7P5XrbxsvH+lxjk5Rv5/Bqf+vsOFuCEFS/jFXwYQWDLogOtHZVVFlUm6c5aZzd4HZwv
h55EzhrVZDJYGhQHaIuzgXUz3auoJB40UhaDT9uwg4ScEi98DfY1FhZw5ELAUPa6DqdZnrcgib0G
AyhRKPX6klrEe/d3jPSrv00LzkKMCGwwSdQkiMw04UlV1SfNRcUPpvO4DUL0aXKrsyRbpcN3/2Ff
3o8ibhZp/W46ldxYwkwJ5WbEWwWe7GczCfXXa+q9TmqANtfGiDgsV118Uc7f6aZgA/m2W2b2J5yq
2ZhGpo0HtEoTLssH2ziAZfTo0AD51hY5xpsKvOmFEJokHQvIaWI+eIojhuM8uqRNpwGCFVl9mKys
4w3ZBNv8NeN9S+ulqBQoTDhnlbaeJJWsoAvMSG+YbwBp4gBNxLgy6Ot/c8UdDen6PVD9m38zk45K
qiGO3s3ewKz1XYYnhmY/gmpWQ3kZhk95evGBuNofBE3fsu0BKo5+lBCxYSZNhEDkJcAdP1GxzVCy
gi/ow7r86qEkMm4THdLWjePMAVVm11fFrvGARg4J5zhwDr3K+91eFL5DvFbSEGBjetLMmCwuXcUi
xRRUi9GX9SI2OmL7ZDs+RgSKI3XUim8HaY85mmam8cB97MCfMk6WeB9B1azNKtFoVBiwhtDHoQUO
E54+H+qJLKExF0jZfH2gxYugRULXLoZJzd8zeaSdVEmEDXs69skCAVTlm68nr4MdzNy7jJL7aECo
DWQi+5I4pDUcrXtLGId9y2Y2DBTzaqHykpg9qvufKKVXYEKG5GrVuq6B9a6pUqVaQ+qUQytKEQmt
Rkv+3FxBxqOTwOEwGiL/cscPO6SljOiB2gdNj5qYWvhXv9ztif/iCbQrvzIzgATXtQ1O4iVakRQI
hEqJdmngRKbLfY8eLTibIAta47mjkFr0VYsaoXoST2thfVrmXdPECrOMQFxmpQLdMqdtZ3fjuUB2
t5/b4rOF/ITRYm1XSs8NyfJxvFivM6HjGmHaWqkBwP+DTHdsp5MMPQfvkwwUpuvdVgAspl3Zsgpk
qPFQVx4cD6j5LYrCnVYXBYS8wGUwNcJFcaCbtsy7pEOQHlAadZSWDpPD4TaXPHzmWr0G6TPxwREP
nC3WqUNdaNYR4k/M1o14iO9NZTmv1rwgkLMQOUgfrPyEKlTuM6pevYhHXP85NEJmXc2U+Lc0WzLk
VaHe7zUrymQu2tVb7o70apUvKaebVFYj7Ng4DssjFWXZIAlcDoTOlXk3rUQ/Ices2hHzOLE4QBqL
JqWP2fgd7TKXQW3b2YDKW7Dp/4uFc1W5ASJt33tJR9JYrfx1R5HVHPQZGHif3W0iWlWn8PHYcTJR
NhZ2R26ETSrMeYdJKJM9ol5MObL7fyDEiyUHeKCpCAt8nKLqVApCexUlA+CK27RTEYlHbp4gRn+G
2u4vjE7sflHGP2eb5VRGqfPJT4y5MyphfknjCEcL0Ni+xAoSuaFbfcvK2/D7HQyOk+1NPDVzOVyF
Wp1eNgjfgdbN91V9D/6LlpIAjwj/lFBk5CmztBA6GCvRho4pG5pT0oe1Kndz2NyZlzba5FzLAiZR
Hat8oYz7ODG2tFydpuNHilGcmdBTX3+pEPXfZyHy5I0F9D6638rUVeAdIM9WbK09v011VcXin6wO
1HrPw1RVBf+6pvVuJQlLDbpMqMNsDATgpZMtLD/xDLdsVC3EgIzLfqVm7ukVfF4mSfwoQT2HNtW6
3WT594wH9Pb32ouzE84P7Pd108Z5+ZdDvxsQVopA+4+vw6y89rSzFJ0IZRVB3/JiCH8GaGI4M6JK
v5QV+ZaLYVX6+o14EaKLjYnuB4mjkK+HTIjmd3+yWn73F3RzhURITd5RkI6QaizX3FsyDfcatrQ6
r2gvSXmGceU5Kg+FxNNglhQB6AWllgSnYfRdB8UUiUyJOO3gtIGvauG8d3FiFk80kcndJJSdFw1k
ZHmzvNDhhv5ACTufcb3lqYu8gLyhwWn4nZHsAlbH5scygR2daoMlhhmdJM2dtUV08hro0xlrDgPr
MxC/7TbRmBVEJnaXhxbB8CVMq/xYnqlH32stpmIM8BgJWjUz0X098XafZjjJIlIbtRgQo9ONGP89
s84VEv7hLasUrjd2y5bY2+koyWNQuBf4qEO50dzLLebGXmCRF4D7MTAqelrMNa2PiGhhqiuiZ9Px
mwvJD3CQXeyArssIaJAhixYjUpiyqvWaP3+zh3x+UCaTx7aaJ257129AChNethhCsy8jB0BJuBUn
1rL+KEr9sBOedeo39/KZSx4U5NA54XUlOWmd9fb5MuP9HBS/pwRQT/8gpM8Zxm9P0n3StGRYoM9f
USZQNhG9MD3VhYAoNRgP6cPtrOOpR6ivg/nnF09lLXVCx9TkY1eiZvGt0L0CjSrr6VKrLxzrZw1E
2SxlWK3a3EJIBi0V1KTa6UOnLImTV8kyYgKWWreJHmc3elN+HUiW7nwphsywAF+dLNc7st79P/Vn
gs49G8PBoi12NO4eCZwbQ7JA12zLcPUN6yDcIze7QEjUV3YzZ9b9EJWwEGhCpaiRqkPgkLb27kjA
eaTx9teL+Qq2sNxM+7n1ETdWKHFmR+QuoV32jJYLxdD31e+BQhNoMbztDqD27chhhP7AQKGugCDP
5tirIXsYQ/N4RQL3Q8zhQ/8GlFy0WlPw5+JK3OGCh56EkRXtIjDmNacY4VvNnCnQLKDGCGuxBaKl
c6hIJTMtrrgYleYD/mU/7WiImFST5iTwDc3dCTVJKULtePOrDa0aETA1n+5sROwBDKNwasBjyCWc
vKqdULTl3xq4X1PzPH2/K/Tc/IEgWaZmcjLDuywrMG3NPHpGpjlBIIMT0GS1+0nn4YhPleUV1vrL
p0MlZYVjN7T/3vycHWwuCmRV3jOrwfSWE2RGGaJc8wR2vN0djR2hgEYZCTuCdFB76VA90Rpzzr9p
p9837vH4i/PPHsP5xSH4ooda6TNOt03tReCNzqYxdUnxo83q1ZevDZ5AYOoB/c12vc8z1E4Vq7od
Dz+TVT2s59eAhWl3s8RxuriuJYZ8SWWPu0lP3toOjUD1/FPHQ3CJMpJETGokiOa2jAbmNk/f7ah8
CVMEHAOFWhcye9yGqETuVcP9hPr8jU9cooTvGEHdrUJVPKeg9dGxJCam1wZ+39E9Fbuzd0HBjpB4
TSQiwanufK8msJnIq9pzoVglH1rvBswNhrgJ6tXC2WOAuHUWcTBVZ6nLMXC6iMUSs7zDHPMEWe3U
hi0kysdWU/QfDZjHZmxs20QsbEUY1l6s/31iq+QeOx34Bj91XqZzRtqWmnMjlvArInpvxdezeE5S
5aEukx2BuUubtPMIHR3eamksCI2Uv0+GBW+HXk3NjTXNGK/EHXq3o+YYTaS5a+06WQCrZ3uUAu0J
FabMa/1Mam9ZPUCxIkA4MWmqvLz87iUwEFIZ7yn9zlU+ofEp4B0E2Qt7ofwK95c9PL8q+1+OxHrq
PN4k+5jJjdpe3iimQIy92ORaz27+ekxKV5bAd1zgg183vnRXzfPnW6YZ6Us0EX43R6/oQkqDrAFo
vbo3111gJDBl4p5vmoygf7K6YURIpXcMG3Mo41BmoZrYwkW4HEi8i1LtMho3HFKMIsfLi4mnwMwc
iMbMJ5garsqcNhbrqbStSaoNOzWVOsUD9oU8BWzcUxm/mARqqI8BP2S8cvrwyEt4NigtTdtpSDZ/
MJqdI2EfrG77aetz7KE6qsOqW2qgnxkP9w1ME5WEHglfJsjyaVm5SFg/cPwT5jo4GkMqdr98ukwC
C8MX2/LshxpDLzz+b/4NQEu7GWbn30H5THpAhbBW8YerbflDvbWOwIwqErC7AsctF2BJD1DruaKT
13FmtOdk7aC03Vhc4dmT27TFl7Rva+DNyDSqQQQ7aEEOuNSg5YJNTg9dFhsJNvX+/gfCe3dcGT5z
gKs0lCjftv5ymVh2tswSmfm139+eGr0xEe7yQ+M4gfTgGNPSI1AvOTze278vv1pfEk0xJUSyy6Mo
TFDCj1p7jyUBgWBRhOJFU5PWsfdqlnI5n8+MdjIRuhB6spDyJuau7QgLbeqN1KroEtSloD+1aFNZ
RxLpQOpL2Q8gAz84SLsfnQAr4yF7s9KBdxxR0nT6B69zJwtMo00kf/JFr+iY3Vlxc0v2SLBnKsCA
P1QqDH6nnCkkewXgJaU64OQuSPPJK7a7duQjDWt0rpe+MkaLAh6b2Brg+v3yNgLy1UH7b8b/k7ua
tSgu1vQluRcqP1in72ZeK2ieS74BqRZk3wSPzhC4m/R1fuuuEvlqLU+76PVYEJDLgr6IOisSVh0I
5P6WdCNQMVt11C7PSZ2ZNMFp+RJrk5y0MODPKgkcD3lZGxi6Pbumas7KHQOszNx8JDp+qveYVMfa
9n0FKEBsIE5CHMHxfx2RCE6+s795aJzNc1eEC/9mfneKhGSBvuVUBf6JcTs+ZPm0uTcfbHH9v6A2
7T5tA+Jnuiv1Di/dfgoAZ2/Ss0rNVTeA3M39+tFSwjDGSrE0CW8trEaKUk4O8NcixTlW1XwfJfg+
2EdISRJEMxC6nncFCNwoE/po9cU+LezrSNb+9ze4M3mPpJlGVdMcueQ9KBzlZzob5hFg985Q71VX
/0lsaCVx9xB9ggyA8rpIw/e3bKxi7K3pdUGupwbaRuJdQqCnxBKKL7OSIouzcUCox86wf7rA6R9S
0vscAX5E/lYS8yYKSnqf/LWMGXqz8pg6DnPn2PZo9EVQIJqnlrvw/wyv+GzgwywY8PgZ5jflFCV6
moanwDTTCb61TC8a5Cf2ukC2RY2xCmYWIUx8uYvoWg9UA8sM9uurXyS5wFGhDls62NCQ7Mot1Av3
W1n4ES+bn/nVv7rCKSfAR3KXnLk5+5fCXdZ669TEK5llCCCqBfB+ojCzbLeiuDgVzHmPTihMu2GP
0a/EAtGoJAL7wYYdFPG/3DH40Tg0xBstZoCywYDl30rPqPCel9yES0JV4q2mTn+LeuDGCLp9YwVn
n03fsl/NiP+9KkYCaGR/B+KdFujXnDMHVfi2bsIithPbsVAktCFR/FgkrRwiPCtA6+jpz46K8sOP
Q9y41iMwjlU7NT8Qx63hc7uiNLFlIuq9T5XpFya0dGJ39Vg6dDCS4yWufBC2APx7x170PRZIirDm
UAjZlJc7ub6mHYjV/hDe1CMTeiOZS8jeIQdY0k76eWT33tkUlJ9g0X2s/Q6shUVZXLTFS3aUsQ9+
JhD7AbpBDiSGMDBFKo/OYXCmGJVgNol9KjjNJm6MieGkqhNhSbK0NY1yAnUDgUqRckKxjaQAW1ju
cuWrFmO/3zNudMjvKY4Y6d/ek79X6ZwOkdTi4TZ5rW+b+wRmUZfE/275ShANfXM8yteFK2S0enYI
bEbmpCcizpwtPnitC6NcIDfhHdPGSNf28oETMeFkT5VFc2BCzRMqMJxPaf365+10wJIAvfu9duV+
ijF7i7dxiy4PVT4QcGUPYTUlNObA2GaBRcjxrHzr84RLoc6CKNo2SF8RIILvlBaU8e0Hs+SWW+zy
FkL6lNWhiTXDWfvsXB730yW9py4ItvmHicF/KL20MuhrBwVdXrVsOFJ88VzJ/0BqUcZigxERPl4l
HlMaWvQRUOXaFZEm2SW/1unAIvFPTd5g7g+ZprLSf3MdLim16Xv7+gDwUM0G5f2Gu9N85fA3gZnw
L0tkH/z4iEt1dvIYrG9vuuAisBhwB3ZY8I3EOnEM9bz7ALpiISs1bVh+qSta9sd8JK0n3AFbDfJv
BCoAqDFodHgBzC4vIUP2Q/kiLT5P9Wa804b6+dzrJ+SxDBbPbtFSUcedcg8W8WuRbNOroyQUPpMg
VcXWIWzN4llmmQ3WGPk+m+n/d5XqOX0pJOc9pA/3HaIUZiqJkFaORhHB7k8v8qBLsPLyZB4MxcK8
L4atxajYfChg+3WQ/lhzbuG5GZXUWUeh0LBDK7KBzPYrZBNB9UqsNAIKvzk93hQA/U1nrYeeKsTz
5aunREsZxAwSU1xLn7aDTdHvOjzHgbAkaO7uNAHCuQoI6rHbjgqiW63Kno8MLn6FSgk9Q0iIrznn
NdbqLkJTYwPldbnCSS/xSa7gwRfM16HhkL1sxbMujUa2G3CBU802BQzv6iaE8IZKdI3k5uXeTgAf
iuv5juaAXeCmZOFCDKqBtqpUdj40QNabE1tTd079r2tGxPNyU2T2DG/sg+42qjAk5xf5emTSZWT+
lae7rT0Ql3PK+8/Jv9qhL4K5rBN6Ndg860jrehljRW+9LyQ0Qq1BG6i8fscdFwk7uShNqUgdeOZG
5gaXd/B8ruHyIt3pfxUWsm2pGCqAnGv1ZAkqkoIKcp2kws0fC5Gxv58VAEtxwnHliq1l+UllSMFe
oGBojwLPledVrpZW72H3FMvZlE1CPY8QyBUe9IB8rzZ+LtFMvVrCd8f2TkPTfT5K25Pq45eIwfxE
UQBu4tW68xhPYoKsTLVGwu0evLN3g7a1ebFqSftYwNht8slF95AxN7t2qGaknigHBLBU5uBGXfil
MJI2ABwitMpjjI1Eju0QwaFr5ZDxJOUIXnnNH0CwKzGXtjtt9X9tmUPw/rttY115GuwsDWCs5Vmm
sJ2hk1MTL1yGYbwR7+dZF6M7Se7yVjfDHcaNk/yj7y8pTRqy3HEax2kVmCf5US7mWR1Ap86XMs3Y
zeXT47gBls5b2fGwTxOKzPWNz7t2rGN5e6r3dz6OkdoYpB5NlDvIpJIDt33nIIvvlqkdE3m8KBwC
xf7H74Ad8mOpeCh4dLkzaPDqJYZYohFisYp/fmw1Ww38diXmz7K36LxTfoOZrJYLu8GhIKAolBVO
rWrVjO6qcI6F/yMWmsBzx2wBizVBJ/iTSQg5zQsNgn19iMxzlzdgQ7OEN+B7UlF+6N+yZMfozYk/
1RBooKpk61sPy7Zp03iMXEjw0Lu+NdeGwwpyF5R0cPI6LOOfyEX7JbAQIjyQSGyOl+RKHbPQOtCW
xKVH/a34FsblSoISiSPc1lBL9YVfkS7Yt7Pa2PU2oF87ygEXNyKf0aBUPuPKZNkp4kVouNnIjtO2
DzSkeuhWwh1AuSOXQ4u52XH0eu04+FQPLihVS/9hk2dpHWg2AZiY32HSirjR8ObfmcD8bPXV8lzD
bxrE+e9zP+qy2II3pUmQQUyPs0VUJmkRvCb+Y8MOEKPHicx+3NA2f2CvHI3MHrWKZMa4PoO9PVhi
qisgGgBjEt1prnJrUTO11DkxS2ofEru3nyVKhIJlk7ZOIB9CujcbrzT+Nb1NwOex2oTG0FLlfFKn
dtwADxC07UMsf3buZ74DtDjPi6wMmQxAt4OpbQP5GFOb6grh9yo0cc2Lyq1UOwKLvOFVcO6/2IPz
pqTr+5Sz667h5uQ8nfD4SsGPQwBne8GFYBnCL/lE4jMaUXkjtPAYRklYTQg0Z9eL8GU7Mv4oojVV
NftxD6vjsoG0GzsDlFnP/fxxe9uYJPBJ5cCz1dzlpaxENhJgrTOBbfCrV5vWthA4YXaBEsT/CiG4
reV9hSCog4rXc9/XpHrCCr0O49hmcSPUPzkcUAN9T1JJJxVZ1U048DS22kCSjBdvBVOsQS20f9MH
asjfW9vYpE4QhlOwsyO7s39yBUztnQKbiKHBjuHshcKKl8D10IEUJubRrOoePhJfh3gjzZcO+bxs
IkhOqpbfdkgkVmtStLDTiwocubCfzn0YY28VpLeXDJP0yu5wY5CM4UU8tMshMH/pbqHdBP2brt/7
Rk68eNaaUUB/rfajCF6wKla+53jpkjMsrq2XvSDJALE7tXPLQOQLp1dtN7V40zvk9ApfBL8V2rYC
vAi40u0HJFRR0tMHTsP67n5KmAc/UmZfr2DbyUP+hW5mSaitBZ1Gkg8uUhbabr0qaxqa30KTnr1c
G1f9mn/w8EWaSTSGipIs8ViNXFSUHZycXZjFWHvmVZEvDy4tlYHJjXtQgBEdrfBRTczEq9jJ5id5
glaCzYTZWY6/5ppotMvlsq74dalk6ye7oSJ5iUwX+xGm5FQAzx6bdZQO4AG+mc1rHM3KauzqxeuJ
a6+X9F1LhezgC6Mq5egfGlKQjMCo2daOF/hzOg45lZ8QB1SWR+nZX4UE2XfciA+io2QCZFTcOQxe
M4TOeHtDhGF8YSpU51Yny8pfiLeOmYpwS0tANHgGrL2Ef8jyiihLw4626NFebPKzUuCo/NxvlCUu
0iZtk/QiTrgbBGoqd5zYDQslnlZQW0m1Azjk3wwWd7YmznTTD2lV2ijpVDMmI/ic60BPvPEcjbhM
CvPV68UDMZ4m0w83xA/wNiAU+lICqbYYyhqoP4Hys2D6bLY4EjJ64RyjpljCgi19joPtoSib1KIf
fPzvugXQ2kKrfqG1bUwa4aXAT4CWUg9eXF17kZzmAWOYMiAev5iARmkTIcs6QnJFkYKja82COGgh
095NaT8TbsNGwjE3WWVROWJZ9XEYuxYZaSHQ5EKOOu6i9JJcgN7sNujg5YoN0Ew2jf5/O7sCCrzU
UbeCW9zQScPDo7T5Vw0E+Cn+fEWL20MoyFn+yYMyJSP82pnrxkuHBX993fsR1yBUb5ypocwjsSrw
BFA+KAOU2YJwquAS7vHNQqcmjyhDwAoleCb07bDAt6jy/U2r07DvB7xCy01v5AaligZesHfSRi7S
pZlG4UG4ORMb8INtdqFK/Wv0r7RoSZEXFaurA5IXH/WGgsM0ca8xkmrG3FkrV9Yo2rdzHkN8AFzM
hr/aalyVHe6wsBIBgRqiyRrkZutWUbX1dvoleA+UwZS15ZKAiAvhMZHkJ5Z3suc8Be+1ts7vJz1d
yB/q+D62tnJoLJc2Icd9sApWDQ==
`protect end_protected
