-- (C) 2001-2022 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 22.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0RKQNHUuNVssiQBbZU64eF/9xIahmrmFx5bQZaB+b4qqqZKaCMF1GYj3RxhKAFrfhrod7pDq4QRW
m/44u2CnrcU0zh2HOnUuMd0bUB0i/TEbteCu1vW/jIMiBYqu6UA79reskr6uhYHud/QUquJ2gtO/
fDyJ58tJZZEnd8YWUNF324sI7tTuEYP8qv+hQNjVm1AXXI70WYHlj3Q4VAFhinghlU0k33bUywGu
x/8i77RX9HrS6zSYP8KDjmKuC+uRWGgP3y9aZgTJuolGgbt0tktqSqNEsaCBsv/8FsOtUtlqNa2q
pcRNiK9ZU/jQ04xciyympgcPN0LoJCWChqb8EQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
4A8QCjCqx6HB0EpzPR58esPDq9TMyEcsm0ollROlmgHts90aDQxeEM3T5w8aSG2FEsSetU4Gfyp4
fWKBlsOhEzgFNGIWIzFwfGtkRyq7ib3jVqGF3jioxpqBXnnFYiO6wqJp0gaD5QN78RpRrrL8EV4W
gX0DGKm8s2J4G30QGyZlaKSensKBgPrvgM6LQEvY54Jw47qr5o7pOY7p3RbduMJWoa+cZWCa4egu
RatjEhqWJElqdJU6l83g4+YzU5Ds6tiRBwWBu+igxC6NaJEnY79q+Cl/hpQJ3In0cLPM7rHoUHf2
sCmXVTReOducqBwD06JZEDafSSaH2s2jujDweqK/lTjvvYvg8mTmhAeNxp/wbHDBLfvLbRzlfTqN
bCRwhIKOzuymMAkhnjRDLeF90Z1oYajSdumV9Nkj9+xE6NkKigIYR7LGd5iPFm4NrTtqRnIyS5cX
oQOC+U+LGt4TdbgxSNtgcDd/ATSwvdQuAP8e+fWOYjbH8sDvg9nGdNYNvpLiszn3dXDUcgz6xzAW
rQ/b8QZogEyrH08CY4Ps3gaJIGCbSxI3/yWMB9V0ZXjJPslkQhP+8n+LuyWV50ItrtBWXEKpqzmY
uY51BedqVCXa1toUwhexre9nGmaNfIZEHhAtXvQPDCvWGu072YXbYefX5cc3XRuwMMQQoX5nlX7b
O0tu4eXMwIAkQ9qLpalODhv0Kl+JjgdwyPe/OZ/yOckLSw7RIzXEQLwEG1rIbHKHDpxZuruShjqO
3glvcwScPqPxlUWUklqWIDtXXL6prM9krLNooNcpxayvQVbqMXe+7ggGW8NRcTe176llKBt9Me/l
Ft3N7IT/7LcId8vAyiJZmej3wQtyn/2vj3bOt5BkJQcZVClnlY4XJcLE+7e6HSx/khNB2hrJnfGc
l/KzV1W5oeH0YlJ6TOKkNeqApHl5jxV/NCYlley/EZYrMoHiO41BmUifiWG4LIoGQEcxggfIXxpj
GJGkU1NEeWaFlQY9Qsq55/Ldp8+xVZTYtkLcBPb46k6GAlKLecjmPDK/kg7WASxHqDCrN5Z4dASU
evUVNOJKz0JydO0L8GMIP+SgUb/F/vklmnhXHfj6yIlvgLeLVSgu/Frjf4On/DfLShsDnJROGc1s
4yVbtAKXvBeC6rblFAVDyFAXegPt7xoFpIzYues/CUkos4wZakNZXPsvUjivlFS5x48cC+X2wo5y
mZ35tsR5H+e8YLIrVUgG0qEzYhp85GPGH3v8I/V+ACOGHuw6tjkVfiqV2TAB6g+ZYNGoxWEkN7Iu
aNIJADoBH63KVY2DazFfyFzAA1k3iEsFC+656Fv9iOfIi0wGdZ9KGfDJ5CvMeRNHmWDtrjYwQOO6
I6m8nQvyxpZ6KGVCW5SY++rL6srqiLrBTNgDpsipw/XmXru7OkBt4vtOTOpWweMqn8cI+GYGFach
cZLhr/sxV8jCqWtuP7lIlcms+Ww5cC90pqbyB5OP5IFu6MjHRDGZXsvirKnRg0xWI9fx7PqYYouh
5nInrqaHs96U94lr1CyqyYMeM/AE7J2CxcJuneKDkVCyuY6xQ8hMbP7ipN3/s30mZHQDqs6lzDKl
LUMivvuTmFfGNdiVVVz322QbJ0NKK7nOQjzRhourVJ3xsfDZey9l/qr9s/PPS+rk6fZRY1SxyGVT
pKa+ReQ3w3UPE7ZSKWBkgBi3+6/jgZva+n4PzjGKC5Wiw4A+TlRvkdEzuFW9uWpLcJb6WPMbxyBx
456kxwH7o2v42Wh6IUN3YzyKJQPUOdYMMAOKiws2Sl5304jsF2HXC2priIVdqbvqqJD8ACElmAu5
Tq/DG78imbSnAP1sy7m2ZsMWz/S/OEXqDv03usC1eYN1cx5Qw0kd/NHw8j54FHPDq8acoBmYMt37
gtKTN78yZO5cgNbIYBOf7rYoJLQtPKJ/7+nuoKBM+JPBxgHwWmDUTC6wdLnQ/jXjo0s1mU8M+Mo7
K39hKUbovV+z7bG+ib+RDIMNAdsT9MygV9864H7+S+8G5Z73fx1TgttATxnh10x8pjBaK0D9SEII
eWCvZ8iwrQxgkjnBjh0vDU0U0ic2751bCrB4KXzE00uEFhwW+lOMedY7YfHs4ruRkcYMfTIBT2ED
KZtQq5X6bg2G/K8BOH4GhBNEQtnMCNgAk/1yUwRY3/o+opUcTtfQ22lGl17Fyn+/qIZ7CZrSEkdN
jHDPUUOixf/awL1ZvQtbq1Hoe6Ms4MG089NUF78M7Swt5AAvhd2adOQNjqesdiExFc0IzARPobmO
DmaDd9TekKVhnsIaTB7wUKK40n3gnhT8Gk1w72MdrDpR+aSW6XcNf+D+dUJzlYXieYjRs/yVAvE4
9V92qqZ1tMlQmPzy2kCK00Nub5l9l7xQ2vS7s2lUGHLbS75LpZ3MPFYCQ3xuC1ZUg/OhGnsXP0Jg
0dGt9kjIkG4DkPv6OWFsouCRid350JJiNSlDrtYaIm6p08Bbg1KDZFn49mDkbMUdX8/unVgeqCWQ
Mvqxpm0CKq83RGWwjBUwC65hozexuMqKTZ3v+rKkQgSAG0G2T+m7c895JCxGSlYssVsxdqjIwlY8
EMB2v9Ac7Xz9vFv58SFJ0GxUoGcAVlp99KtzQfV7wPsdpPsZPkjBbTzbqTjOf2OrvS1S7epvXM2x
NvCEKE8dSOi+ZeUFTwHiku3CJCZP9Hszld4bpiGyaQ1w/tDS3Xsmg3ACIp2I//MIZiSB629/BX3w
sXOIZrNe5iqMKD6zs0+SL8i5Zul99u+o3SknnnUMzKQ2Lc1rPNxI9+0uxXplwTkI+iW63LQGX5Rn
U9TVkO8R21pHVff1jXw6ZFAwZjl4uJL9Zzq1cF7Hl8w2MWhEuiZjQ9WG7ZyKH2DazFml1RrR1m+P
MzClC9yhBxWf12pG2/VXlQ2oQGb88MuJlPMxopUpxfg0bSjiE8TuEvZm/3vDLSQTtrMwrBknaB1x
wdH5c78L2A0ilpcN7tIJ6EZNT4BiXJqf8Y52hYD+97oHipj8+0i96FHqE5V/j1V0xIKEMNJjMzj5
eOkczgKMK80E1Snp4yGj71gFRw/bjPqGkXfeWy+4wSeSVsEeT8sUJxfjpx+OPlPZN7iY42OdN23v
a005/uU+GjoB8eH5ZIJice6gxvU1nB0X2LyqLKYyOfdVDLTJEJXxWcsC8Iyb8HoyNloMkjPyZnPo
cYyQVIpY8/7ILRRvFXI0BuA1hrimFM3BLZhDVWRSWprWDx3WK7bvRIxNG/dh9B4DeSWZ4rAwi84U
bFQq0mzrHZ/+2z6CRQ6sAn0LGdbRfnxd1CUSKQERcRYUK+PAQre1c6owUEMupN0mtCbccLrlFntz
cLOZgY8P1z0zkEWVgc0KRCAUhBpP0+hCezgc36ZCdEBtGDBvbnvkfkqCpycx4kgQGuR8IZ1EP9G0
WEsUJNnjTApzU04ynAM3FEP9K5ZndWWh6MEihAB+Ucbtv3OOoEUYNuCEuNS9TR3z0fwdkIvPJHH+
6rgYxzV9UQUU+MAmvGUh1wg1X4+cH59fkqtyXBxm/Hk8U9sBtpUlT+6fanZxcAB25JmMDuWfuW0D
rapLH/GJFN0K6k4UXdt3d4WxYiVv/CPQToL6rfwg0BUZAW+t6WN4nMqPIr5G5O0nWIerGu4gUM1a
wuCmaV5uFOqF6dJJWkKwL2YQBpTpeI0SaD3um+b8t06wzrqgToDl5Wx4b8MDjBN/XcEu3gmfAP2J
o3pzLbauivPVp1sqtkupbKg2Wpbqokkle5BkpbE+Rec2O9UXh+K74sPxsUAuMyaXkq9Wz2BVIqsi
4a3VpGCTOMXqQyOkzrbOk7Iq4LDt9uOS6EPxIl2MAclFzXCNkBIxMmQyUYlivrDJ4QiynJH9xUc+
koWkjcCpYIQ9QHlosPYlMr0/nSc/bwEtIl/KVcSLuR3H8zv59CCZbCUXw15NPMwtY64Hi473nTfB
nXVjDQmK07M7/lvmekCIsl23HZFJq00Yyj5sivZUxYUbOhAMQPfE0gpoEGSjP9+lntP4cb7BZvzg
VtVqUXRAuBENeqXfEA8lwytoXoF2DniYxxZ/CUTmRfQN1sHCPRv279WNa5kvhzDg+aDJy4hdNLRz
ufHS+kEnMIl76JYx7Rd+0VQUZ5zJGqY6dfD9mC9BMrZl3E8+qiM1T2rdR8AhueZwCL8fq2vCKfxr
5qY2Iiya7d7ylqn07e8F97JhhiFZ2NdpN+BldmFaLRtfOI4KPfs/jYSMCaZdwXWYLt6UhV9wgnuL
WOX4SoRXsA0d7hBd2QCw9GdazWEVgZ1PlhuftqH6NE7w3sz6AWcNnj9WOsXhyNLnmOudqUEl3aNR
tAmROvMiZzkKmoFjn7aZCXLCJVC3d/iQ8GmPJj8l5oTxnZAEMRmSg1w3bl/DSawYqoVHPU15yyfY
9gXYrLYhqA5ov0rPonXejd1EkvamWA9dFHyii3mOVfbkswJJ30HhsmoV54xM6TxBEjHtgqIfEKK0
6C3JRhX/l61pBuOPFAIAVuFq/TmlTPdvSTTMMjrczOX+r5S7gAZevSvC9gq41yuPp+CxKQzt3Rww
Ait7T3P2j+TtHit4seBa+f7pn2yr0q1OKheCt3qAhsNwcwM54r63p9azYGNMLxeN3WZ5geZdDOjb
qYmSxorcf6iuAqroBLivhwwlnic40/KvGpZG37Gzidoi1Beq10DGYIlzSYybqs9ka55a6yfaGXp2
mjqju8lovGzh5oRKhlknc6jXpPXxQH1xUiKN5csA5V51ziXthaamW9HM0KLhvJr34zGxLQF0k4QT
tHHyL7lrBKAtG8eJufAfdiRPNAty9Bn0PKssuPsFbwh4r4RsIIZ5STV9JOmgorCNF4LtMKbAQ2IK
dJ55htPskg3R3D6Bo3D9DF3uB4TgEaQHgKFZbbzfoKtydRgDWj6vShu/8/1+Ybl0RS4JVLug15eV
rMk8DaYDc3/weNNmqbnjIWGDU3EgioIGs7lO3IsyEF7NMLjCxN5AqJ/PoxU+nZVXvxTfbO9VQJ/Z
DBbvCC8u1YMSkHcYxFgzERe9aq/s4YeSoOGyS9OGuCKaewGlwOu/FOaYtetNmIaGMUWDD1O+IZTR
6Lzs8kpVXHLRTGXw3gtrCz2HZA3qW+7kKZ83SrVWVhFBPKRpJQlvK4RD5GZ6bxppk0HIxm4OiHgo
qPoY76VXdQeei1DoXzzkeXQanEpThENWvAqZ9GljLNKjKuW2p+XVEjsx6tckgKV/GHiNh11huMA2
jCg0pW6WGgSeMXE7kzihfNUeU0KZC7l7tS9215PwSc2eX0b8GomjesT8NAYT0sRyp1opBfK8mIpp
qdz6b6DCufDZuNH8wi8P7uV9JGb6IcSRNTwkIKpGWpJBHBLbtEEZgUa9FB/iMSM+kXTf0qqftnMS
IyY93SSV0wwgg1pCwgye5W+wTAdcufA6TJKbfb9Shj26XO++tWvopODyr1JeR5QY1ylh+tGWDGmN
H9hYbX3ekMdWtSpmcZyBcFCCPFB1cjBj1W3rac0GLhhxmdFNKI35NKoTrbzQNYv/iyVw/e485QhW
iHeK0HDrIJuJGIJ+xwLjZDyepwyPP/n40eKwJ85bzfnj+DTHgp83NdEazFwmhtVEMx/Ek37cbYVn
oagCiyv/Im3rp82t2N/CkZwF9Imgw0HmUWmb9YcrO+zbWiJG+WkJ9VUDh6z3BLQ2pC2FBVT43dgi
BDevB9yQuR7fVpHBuvB26RD/gAcOxx7paCwj7Zxvbw25rkttOJp0FP7hroKO+HBkwzvMYgiI8Iyr
pTXLsCQ7AS9GLvyDPpBrd0P86Tyga1OS44qtPPLOyWN9OxyngqdbmYwuMFDh6/kBevEuDGNEZBXs
V2Q7tP7oeYJU1aAVBjvj+oiJEcwOjPQ13cuZLshmlBYepxQ5ir0dx6yK8ACMucTNPL0ZFDkKZ4K3
PpazR5BIDpOvuh3RoebpDivsJku1vh+IqRVLnqJJlnC0p3PWKYLM3Ig4K7xhg4z6ZwUfULqWKDb3
zF89/0FLrY4VbnALHpDyHKKuFQAL6TnGOo9tUgTdzMJ9VNX8qqdouK3MKMoT+NVz/weVKxh5Kl1K
J2xJMtjQYC716mUcoGPe5PCK7wThqQsmDYqvvNxHYsg0tnaBEPZNwuk+RkA49S+1CBkpMxkAUxCR
L/K4a9ENHB3DH58YQm0HhFoTEsBfwxMzVG5UnnQ++qtBySVDVNDBhhXc8sU8jeW3uiiqBKbfZhyp
r55declUcNth5SADvLvLFhOUchc/F+45/v1QXDRKuPoUR5ruRMA4P4Q0CsDiIZX0uanfaFnH4EUf
ra1xMHzTQOF+IvU4KpmnG+gBjJMgEPj22XWFXOS+ew5V6s/5xM3hn2QgMrGuUPVOhNefEkkJ6RUY
2OMgXhjtCK4vgRN3SyY7sYTLQVYMQWe+G3u9KGUPaE5uFiFFAq/9bdjSJGBfBHdUARDuDq/DtBit
dyaq+QutXyZFkXI+cjYEBVEnjiCSMlmQUUfl6Do3UlYwjPo5k5VWtq9adppQNzfkatMlDY3o69k3
axb8F3Vhm0ceaJaIKND5lSDcOkQ6L/d/dKnjp2XY2nCKYrNjkazj87Wq8HX92TrE4NvF0TZMN2m3
/cKqJL9JDC9g8IMB0Rns3bj+LiPHeSv1V40wAgbAcWzBH3mg00F5VedH3ibTf79kHKZ1ENVEHV36
zzD3zX5/7kuGjyda8xks2LdTSuHili9n4PUxHm+ej5ChIQQn5rZVruyTrQ7xJ0DRtP4NshmXjFgQ
q0AdoLJNJemfvNvGN9i+EFtUfCB8r8wwTFtCdJaSE/amgidBzkiimh4HEEIyuNZUDb/skas521XL
7RB4aJhm6xhQcyx1avQVQfrrVoAsedEXAtEfYde89KEb8YZQj9YbG8Rj+nn0YRoE3dNJigV7/bKy
FjM/MhG0ySNaNhX2XKr3CTs2gHi0ZXq8fRWpjFsya1YZ8GBQKpxzGpJqjqRJ2EDB+yHHVBOvuSsy
LqTDOXnqQLovjnOD+MZjDK0fLfNa6Ih0bNX6nKi4ujJjWjOcqYZeieMcUVGLuSERfP17XB6SeuHM
Yzu11pPuuKwfSLhc7gUyYRDEKjQ55Gblx0i2jFqJFlOEFxkK3B2aaz0e1Uei8MFJWwVOcdMTUE9I
0qaYh5u/fy15YlZCDpBCsSfT8FMcQTxI5nmVC0J3w7NtXpoRN+PQZVb0+uwmLjeyXp92Z/XHK3Oa
Zbwu3zfZmaWKkO//hZlsRTgEojkpKkPnAz83kUzPZCjcp0SRZuwCn/O6daBBi6SeMMGZp5yKWoDN
EQ3HjABWozAlp7LW4v8cJ+TmJ7Q6bQrr11UL5qkSw1/k6Lv/RUB0xkFr8u4ZCoS2tO6uCfPtf12v
lLHDf7rMnCmomM4fxFCGxcFlJmpAduR53KrFMpk2kpyCj2dQN5pQwPtKfFCASLUjyuRKxU8zVF7B
VPE4PouU1svY+Pr3rg+D1IU6Lb8m4McASCTgZR0wPd9C9owwYNznc8Si2sFprRRohS2PYVMghNOV
42x5CDO06RJnfo651clZOG+XKullwKB7UeeJppGDZDvav88L1MdpcIRuQIOR4aNjLqdEeKmpZvTt
3kxcPaQ84fYTv0gMPC4Vy8pG+xKNZeWPin/0QJqLXs7GgZ4Mj4KLxwVAdGlRgfenAuJKUxxkE3iU
3Sq7WNzLbD2+XAifxJunmd8X/6Ve2VmaC7zStvtDl9arCRstjEyAQLmeqlW4nf+Vdb8ieS40PxT4
2+DfDQWcIoZHSxcoX8EjnZBIYC+p59ooCNOmFZYKrSrqJuQEfARwf5FDIHGLPEFnbBkUwT3MDmAl
0udU3IEZotTTeZqrlU32YI+Y94vBEf45Mx0P9SmkVjn5DdKShm+kFtdWjng9f+jgA6KD43aV3kuh
Bpt8FTx+sTtPRxDrGfQgSFcLGjpwfy2o0D8OqvXu9LBVzKsoIn6YjSw6XMR15wDfLrwgg3z0Sk5h
jYcXgf0PRXLbh2EceuZ5IVizezKPJh0ycS//W+NKFXi6M3iPA5ucK3nd1f2LBm4l40ialFzY9EPF
lhJrgnUe8iCUh0egnDbGW0dHCHTI3sTZmr6173B3oTYbMknaoFXW27KeZUHyHCSxqv27lAtLA8Bj
e/HdP0kzmg7rurLi5tevpOyJNELwOYeUcxd38555ggzjUYhXDKOWjua+KjOqs3aKKGwBjws0cCzL
c9+oaVsGHOXC9+/MPNf4XSL8S/LHTo2s8hIJ9QwsrL/NEpe5jnUO6SEsN1ScrjxbCPHZMo34rZz3
vxrhqzUnPzCuoZXXMKt0m8jrHjUUFRdRnrGJHEncdkQi47umHHcJTQS+EeIAXuIVNvkyAdJwVBbZ
AaZanUwSe6Q9TJVL59OI6i7QWLMqc/tlNAw0eCVHSriZVp2nqEc8W1YU+IODmNJNvGlIdHBCO79V
/bWpTTqvtk34g7krOd1D8GnWZWSv403iXfxAYTBxKwM1/HhPKb+IVFfi4klh+6cGpLBLffuxIoso
qAysIAiAcOPwSbqoddnWdognnVlUsD+qtX+xfF2XVIgOwuWQqpISZ1h12OxLLpX/GYY1cM3G0ivo
EFHrESXjKUGI3czl94BSBAtFQtg6HrcI+uM/Bx/GjBQowaciml0YNnvzWwwzSRVR7rnTAw4R9qlP
unCg41m+7e+dNrlp64PoM1vESW2VvbubF5YQcpSZUiJ5F2eHcHg1HJsXlbkbv6CDuOSrWDsQZm4t
dcf0SLvFTIzAvGTGXr/BXdAGSlKTG6K23yyI2mzyq/7hH7KkO65voFRQYhP9j+y543xzKxBYxAMx
xoZ1WyLZpYXM1G3LNMd4NATLAc+izTG+QZtnPdw8RijuPrz38lgbtthm7my2TZyVtcXsQMI0Y1M4
GqPhQ0CQpHmEE4Cvj7ncHau8av27e8t7B/uiimOLgHkEPYU1gWpthi+DVMTgcSRTjHEYOiNsn6Bh
jvojwTzWvs4haPKMcdCNM1kr+lJn+u1N7GEfb7pJgOb5qla7Xiw5G49bk1Yp39SkqgUnjJ256bEz
77SKpOlX0owBFX6d4CSl6P7eRmra8VZMDjkQ1b6YLcQ1hbYrIUEHJPsEjLz6x4xB4utb8Q3IoOKk
+kD8oOqQRCdJo7Fa8KMCzPDleY0tz1kJyo1xLBe9Mm2slc6nTzbCe7J26daR4q2YSSVpaTQXst3c
r6Y+iPYGUc5Nnrd/vJXcmLggC34TUnzo4qO0KEfy0d1c4MKy/YHGRH/6mdapVZSl4y655w/5x0JX
RIrfaSnCnfuy+lSOYHfYWVoI4Bu8NJUzVnkfQ761yZTuAdyiYQ2JodKL1TPNcOh7Ul+O1mNGyN3m
aAgE6dbGcDkB315GAeKLzDGo57ONsbx5v0MmR2E/LDuriwfWd6bOklfyGYML4qqJFINDL1Mmqfpe
GVq2wYB26it1VCRI0HP9WTS6rDttw2uhXAdv7LTuv3ft6gEmVz05Ow8cMh7ZT9jT5u0OU8izlkik
eH5zIhqvoSLS/GhdFtIzj3e1S8AOy7asd4ytsXMRDR0+w2dBHNzrSFxtUgz9CS6GPjW/1EIaxHr6
8ktTyTiP5v4+3cKz45FRkk7l/qRkCiXU+BCN+fkwJLxPm/7ObNWgzv4UIen0uiLAa96U+Hi6glNz
kpex/PAcWSSJYHu9ZI0jJYeazFai6i1bKnzNeevooWGSuFlKRjWP4DquWcjmZfFO+lsOcBdY5jUW
m4fhFWSEuDzhJazYoBzOdtEscKvySUBHPlufpHb0/FkekPmXnK6qADufzsIK9a7gcFBywlobw8hz
J583fvq8YfA+tDEQz1Sd0VpT8ImIaJE2LL8L4uIVQzHp8C743jPMtnHqGl91dc4LsbgWk2Um4At+
IAQOxYfSipv5qbqcO9q0aVLTls5x+Wgfu+/ob/2k3JWQ2Ur5jFK72GcksmlhPXJGFSAQf9c9W/qF
uc7nuoyyR4ORYrwKNGV/ReJOt/s1lL73GLiFbDwD/kpTQh9QTQyJbXZm7R2fCFH/jKLSMRsaehh4
V7xhQx49xeFt+3+qanPH74w8CJORRsN1MRnBY5mftZwWuKzUsf77OzlDgiwlw5h+xbUP2P9UCHVh
NSAaw6+sKshhMN3H9ccKoj7Ki9G9QhFtPuT3bQIiB4zBS4Hwy4tRhh65Rmix5065BK1Dy0uFUi5c
PUYFpnrI/IBuTn7fTmx2+Ci8OAT/wdfSXhIwU1coPRtoeS9TGN/+DpebrUnJL69eSHoY1Wf+iA5q
ZNo5ErOGBKfyidJ7PapAa25+cFQN20hTPIfzuIAPPU5YOs3WxQnAphjzvLjpB8avlbx8bV7JS6R2
KTjAandNxZfw6EW7RQRaotqlnXj3N5hLglRqpd/KfORslCujHJqJ6rXX3OAviWqmRmUOEa2hgQ1G
cpd4yBZoGJSEKi0jq3EMZmPs43wdA/D/VRsigvsRoLPbhfj3I6QXB0MSmI+jLAXlfZmC7y2oLLg+
68L/53Av1XLacAdyowkD4htkMwh9nTZOjy9suwoJxoL9qycw7RkdfXAZp4zMnQMN4/Z95IMlNBbA
x7Ak4ZdbBWRj7GAIbK9c9Jz9t3WXj/+GCa/DSVELnKG1loDWM+O9mCKkLuBJFO2FUt/MZUUFTb+l
loPNsS4vQAzGQ/tY73+HddopW8L/2JY7FSK+seDrBnDd66vVFtOKqH6+dO+aEsBNnQewBPuBh1ap
o99mHvdAdf3uBppNul0vBUqI+pX2ytuCBmvjHXmbN1u/Yo5Cz6WiL2NBBUyuSW2ikxL0Cj2znIyA
ReQbHKMwmAY3BDiNaHrwfkvs4mTtKoj7gr3SqDjloK+MAvpLRc3yw7jAcwZLOLGjCB3UY6yMVfWN
2bowRuTSSly57eu3sSkJQNBvyu6JtKB4d15PCoDAnePcqqBcmDLDF14EtMyQM4HdiD97qYa1dxlb
yQZhnIEpAtccwNTLhWoDhe1QMnoC/vokHjEKRZQy1UBsWWpGHNoB92NoHpRWODle+7w2DwOSJxUE
gOtgRPOCzzm0wAIStX4f0zA8a+7Rwsd0EttrjfCN/iT8ChcD55pD6KZmc9j6IBVhoDXJngOZ+8mC
kSzQf3kJXdpoNczagJaS26kymfdGV33hKrcFxPbIAIZuPtJ5N6wekYAjcioxIxxVKSl92HOhfSlK
ztm0CwusOgP6JwXMnzCWFBcuEwo5MkE4viUGf0Wd5oUjmVv1bhJ+fes+EWFzTxcfA1jJ/KJS2YPd
dPgWoJEme9ooDa/T0MpX/npiP02q+YY4OXspOhgoIUqyCd/gj89aJ8d1gb9lHqoO0Mqc3NMhY+kx
9xAWD3bnXzzXNxdx0ptoFhJ3OASEI/gBYdM1XYP1Q7k+FYrsllV1nHrLB1VqBJSpgx8st3yrNtlK
DA2TqmCNDsNJNTv5dJB+IXBB702kEacOaI+ZoItwJ4x4xUQwX/Ac4vjmWqKbVtYfdr5aoV8b7NY9
QIYQP5+iLYiuvDpNdsxMVoDeL7BOfT7HaCM4ApiZ6y0JvdDpvGWOHheit5+938ZGeGPVHB3xbm+6
Vaq5U1KJ7MJVVdq4mnpZoc8Q+l5Omwi3sZh++rBs+xhP0br7KOTm7vSnd+olVE5nYF4W8Di96Cf2
THW+NPLP/7FuOHAngMseOS9WHV5+UbLaTadF3Wek29+kjaC7bP2ZIQAlD177loarnLNxpyCnDtJp
+E+e6q9WX3x0KP7AD80iKRfTEA94agNcWaG6YOyqu0OApLa9Vjg6RWDCS8ndQgI9rL3ES+iMq/xa
qjmrUFPhBHJ3jxPYkEF4jdXMxwlEQcJCb3tMl/phIg8l3QuoOII95tsX/gBz+frq+fs8QFuK3Tmk
RxoLm923cDuAkbkf9RjOjdLf+2OvOVO2mY8W4nlSVMQbY4TJz6mXmEolrvlGBaWTgfe6Nsn1tFNO
og6i5yn7eJNwEGs/fs2EH566+0I9FXAGlZImNFqEMPweECM/MCPUBUXA7LRWHuIyN2hhqz4xMPIM
jW2ZnA764NMgZW9y3eiT1si2PVY2yVpeMshGTVDTfkE4L1Idm120jr8zjv5V9zCqdTkhsOTYwEpA
wAbx9OeXZY0GkHXZss5stev7r/02AuVW+LAk9LaQ/haX6dtFcl7YudTVbmmcZI+8N5+YNOsr0+Jh
+Y5iYySJ4dpqXWN9f0fT1Du2PspCCIGrRE3Yz0eyFEtFX+rPJyuqI5ruI1dAL8dgZ5HyTYlP1pai
HOWoZTB32Pwo5CcB1sVLoMRGCfh1pfOsUMDJ6kPNe0LWu3Rta+fGsjp0duGJjFC5+pZdP/ZSUPol
QYDpYwf4XfIBjKAUPFXUS0242oKaUyb/2GVM0ekS7/Ftg+jGU9K7kxHTqBQ+FnNZggJVTM0Hd390
fkm5S2N6SS4/U9nj3II8qGeRKM9q6zkRudNqUveyRtA+qSNopS41FAVY6C69yXgHmTZftQ+0ZG4g
krsb2x0a/w4orcVYSrRUYxZegLVN+CmyyacYK7REQTetjg7CzMOMDc+0UbUYGuOyORnncrsdRA10
V7ew4oTexkkY4TbvDRlHl5vIln7vPnwZC0csYWB6LEQ1MGjlG48bax8oZMijOmIEm7tJXnQSTEgB
ilnkUTfZDqJtV/+eqsU33fKeV/7fjJRyQCSd745iNaRnc8H7lHZzKrk/ANqBCYQgJUVxP9h11syn
YTWv/bg8fPMcWxATJvnWrXd6xBHZk34LLbbEzxBnfiAn2h9h63MgQIUScTOzMi8fqpP0kmJfdypZ
d1Kn79WjG1WJhm02cnGj0GDsdEdwR7FosLxyRq4JbDXMkGTkQY4OsYLV5ca4s3+Zy3ksENgMhN4C
Rm1HlRoGDGSBTmyzsuH+4kQX8J3rl9wxRzY0H51waxHSw8J7IA9GoqrbZGq7aSrftULipDkLk/Tc
27zjBwITXwV5QywG2LiceOM5TUfwu364DZE/KTPxkx1//qrwk4NC1dVnpO4ygPyv6JjjsdOgIyb8
fU8WWMbyW/teDQ+FLFgH+Ju0+8ZFvQXiqQIRrcIiW4QYn+nKB3Q+4BWr1DtKv7vPb1p3jDfqy8/K
JhkBQ/mt48f45uX6be5Creq42IJwVWeFeMcKvaz6oEKIFrqJROZynDlqhyFxwm8imkKFlhKbVr4A
jTdQiHmna+yYq8wGNlxYiEQQLhkbm7Fr1fLBf5lN/2tiaRgHcjVRoeLm9CRFVZKGknxaQDcRMFca
4YFMH93vGaVdG81l6pVTzh5cj1mAt8cdjkQ79ReofUzaT06uW5s+WIuJluzZ6iVbds/AbOp5bFb5
4Bp0yPUKJQWwQSVLrQmOJwQsJv0zkuQO4h7N23R7aoMt+33vi7J1qGp6LCk4pCoKOv/VcD4q/sb4
+9dXypvUsaFz2p66GHWV9DdEKUweIPkAwrV6EF0LQObpUo4OB/4igVG5z2TWnGC4OaMYHzaaqfPR
+swWFGyqKyag2tkc8PEIvPqXjuB9fr9ImxC+tHli6Q93KwetKdJN+s5e6WLNezHQxxFCqx5+wbsd
UfECju7+Hf4Lc8giEEQawlf1wgIxLRMAWcIDEuIW6CreX/c7QH4H7h4QALXAl5VkUtBA+5ey2Gzt
CgdFFDbkpLOE6UNWRKFJsdj09CDvRhm0qlgWl0qLSQKk3AGMG97ofClwfYn9lrggU4hl5ISXeCJB
/nKXcgT3gjga1U2xuEkXUTOArdZ6abMvmJpK6qvRctBWldcL+lSCt+g2KP/694Tzonrd3kFTBvZm
X0VgotnmmrgnRogLJF6p5Pe68jUtmdyqCEkTlqqfK/e9FPn0PmchK2mT3Sq9wh5C5QfIYOv2tNZ2
3B6FxvXYj9kF4g2welRMmfNtsHU1lr3JwTXYrkfUbrOzz/K1r/moWseN1NWUH24aL3hJLba5bmvG
2xDzOKdu2TN/S8vYTG3m4a4LwmOqoZ4mXjdUYO8BjIw7SbBqUlnBMdVZ0YrvVxcT5nV++5d7xbLR
bz374LtG3mRsQ8p8j0/dOxxGqZYj9k0ASInagsKuU/UJtrtiz5MT8orBcQIK421bsHCTOLWsBo0y
XRzf3h91T5x+i0lWoHa5KLta+CuqxjjlJKkVVwW3eHMcwmZt1M2qpCH2BCzMDEOulu1e5dcoWBbm
HOJXb1iRDkrngAW1J8XVGtp8syrXdg6rZHY/YpZUut7kR6xXUUwGsbR5dXSbaC4UoXQowy2+ThWN
Po9LZnzqeC2WmIvvPjatA7Y9cMORjraICpYGJEPGbE6jydbGopAyFQR8iCS4oH+JwVkW6Z9E61Fs
oerdpR2yDqVLE/F/l9pYhpURlVoQIxbfH2mMVXN8n0EJrnWXaKrmCRdnPNdcFpvUH9A41APZ/lTZ
2SJyu5JK/WN8PeKvJQGJCrJUZmwjTnxb5TLROsEo1wF+jgjjGqHREKVP9cfYSsEWW2Iq0lhKePqM
17P8cUsOTY2/OGCiYXm4fRcQmjeVEJxvZXg7R51ZiHocCEHD6gXaR3ou6bZkMV5eOLYFaW9o2/B+
fH31oVL0u/o6eutxX1sJXDp1bVdbZVCSuLJoPVXqC3PYwNLKrHKUEmQkF7edLLET56T3OjVzzH5h
h4jiGdJyDzy65ow/M1hjtkVGSMvUJoCZKHD/KK5/AI0Z58hLFT7zUSZaKF2OoxqlVuJyLfLsMOfH
IdzY8iJjAstZKgTtznzvWk1Ai5w+vNj9m6N+FrZq1zkMn0ca8RUiYcnXOBTomGXYqlus4kiBxPds
zdNKcpM+xSYwdsfuSF/ZAiMqX7WKL0kv5xWVh9ynDr3sO4cHqrxlszem3UX83SEN/s2T5cspQknA
AtJMcAeSsHKpW3trNjUAatPn9X0zN5uwF/zmCaWdOr1jT1BrAOXUJqV1ka1TCNUOoJVrzOv8KZJF
vn9QAh45kKMpFStbjB4MeHgsCdCWRg47ZAPX2bwQnoqGSzEKGneeAUaowyuNrfrn+cMsAXUIhZep
iHJSUZ1y5ykITInQgShStOilih3udyerLlLMhJ7XyfTfnfwX1mEZ3gE3J7HkhPBokOrc9+RN9Qdj
1/vDGOYPxn+95wcPzsvRKt0l8qHYyLQDFZAyC+fOLerxyxlheFP4XKldAewSexSK1HitURrvsAIi
T65GH/EbkJmf7Sg1E5PeHBZEIzGf6bOipa2rbwGccwqwLdA3Wr+X0XlFz6u6eAoeqVLgTBfMy+J6
oO7LqTJ4fmvsHsap4QUXFHv24ZDO3XiwwAXcCPQwc42/qL4hA/bg25AsTAXB1A2YSbCkaR0eVPCK
AyAAUj1feEf7FH3batP0YdmIKWB6cVjOBZKKukfbHztLJjUL3olfUgwcZWCPtW3v01+XLFwj9/a1
YzMAiCVUmHJXZyl2UBn5ptbywnc/oT3rWJZAUB0/g7bBhezTo7AX8TSAlQkw1WcXfsr9KkwV+XSq
UovE0snALUObtg5d41GwG6uayrNWxko2SsokbWNizOfiEmD7Qmg2aX+i7GoGPjn6VfqRXGCsxHw0
z9LHP/wIvXLLfz0o2vi4/w9UhbtXk+YFHzPfsSPFftKKYQDfMMzm3My5ykjq/e3lgVPpXI6d+a0+
8fryxUqYD8xR46mEwP7zNJRifF0+v+VgAFk2iLaT2N6EAuzLfxynUutI9IW3S49LYYTgw9Xzcor6
yU3ow+cEmkjCxkLfrKARtoiy65EEoGyANaEbdhSG4yxouXttsNNsh8cRdsdDtLwjn648nMQkkCIq
smL3qAt8vOVHvxH/a1/cyFoSisuQIlQEw0ybpHY4bvo8z28yK28HkA5JhvFZMrRSvB9DXiF7X8F/
jKfqmpT7ztH8exHxuQq+s9kYNYf6hk9/8a3056NSKEfQqOmDOciEnr6qqwaLuE6Ta5nMUZMjrgU6
K2WCsh4HYToZvaaQM7BzlahbHU9MqSAir8K2SM5Y8L24+tpFstqZsl6g2vmju7oqmTfDEwprDH1n
t6YyuCqkPevtGg9BCHljAyxrj9pBKJaOapwc0eWZi0HsPIXjL7neg3r0lgczEnHarf7td66Xzm0m
+0iFQ3e5MPtGzEx/jcHY+fH05cxRXnjWf2+rjZuWPzjobiCOJQ0Td05p2ZxJoYj0rTGzgIxvgVC/
H86SgKwfKs7QSI2SvEt0ENUhZzyt0jf1fdh9bwr/dvsLAo4YY8GwD05e+NtE0G+SU0gDbjaQhVLD
+3CoT+xesp6WXhBaUdqdEALAOVaoRnyGNFXvys2Ktji3lpxjDuGLDqt8cIo/yn7M4iAxa3ikrgyi
V/9lPCmD5NkiNJcjReEoMXNmVvK4Zh0bq4YoUs3rzwsJ70OD4dGlpnNJ7aub0tuLWC/iWBLCIS/k
iXfGoV4GWkbdJo3rypEqFHZvpsB2lFg4t4jC6Z9qgFAFu6QhCtbqcbw43ODnwzoz3PpMoO+l/iNg
55hUSndDKNgEOfxgY3MuEDHMNRkQFWUtTIMzAd4WN7XsWXolVGTuJkYnJNb4ativiGQRK9QN8lju
WkpTx2gm5V/0IDdPHlRhUXi6U/Cai0uzpT9+14PTKpRJ3DitBABOnQNrijVdTerkunWTQpP4dOWl
yUJhOzj+mN57e9prPDMzu5cT/ytEFNd8t450R7qnIZ9UYLLqeruRAQBHbnXm1L3TWgQ1ww5aLSPK
ikUU/X2w3Zw5T2SVntWMagbLKYfFc7WQMb/KkC2Mb+6mTL2M9/FUVOBxEcEdIjkWY6Jz4ZTfoOH3
IbcA/bfeEORF9Dc4g31EnDaHyX7vYymnPThuecUK6rgPwtRceaetCcPD4+KO1JoDBD9vbuPuQMF0
0iG1Y8sMKQY7NFMebzQbk1AXAN5jq9MlNqDKnyaZKQYPh0iUzHKLLWFG2jMHUJHb7sv6tn+3rh1n
VohFhx47njEGyJVGmUe4/iVxP3D5nv9WnkDqW1MoSoaEiyj+FhYQ2G3r39VH+DdF4xAtBftTOAgB
viknRfQac2dDwXOLHmy+qO1XPwsBPwpPztT1x/ZBJ2lM9M6a0YqpdaY0q+d6bTaik++iL1fpoID2
5PaIEGMKzS+UOt0lS0R4SSoE2Qgbj6oye5j+uwOGqVwbcfie9lEHXXqp06SvTeFKcjKJAvcnJ9yw
AIb8hMznpjMPT3FS2O4dkg1l48JmUelQTpfcVz9Xt4calfWIxBuOHztCwR6TmkflaH/jmiTvJOz2
kT4gKNTScmZvFMerdSqkDKVIIVFDcaZOGIzRhYuc+j/ZXiVvBFxbu24q+sQV/FRmx0QD/BQlpIzO
I0lrDlzX+Xq2RxV3TjE5s5fKe1TkOsdu1BI1SEbGvHNHigg9671rhiPIP/fCqu25MUXe1G8brXpO
JmdWSopzkBhwOsPKOSSoJiIBRUthtNntkBTFCgq4wpDDFHAFfP7BvX3Du2WrNzra5D24bSSOtyRY
FCdsqQUia7OG2njFCareHMFaamXJn6XH5Qsv9Ej0e3eSwKykoaTG04RhcZfYK2ANroFfcmMQDYeJ
Vb52drKF42SLPyi/462NZgPFeuDI85VW7HFyEeuw6BOz2SFwVc+tM9yqJOrhmrwCrH3vn9xco1JQ
g+t8p1EmZevd3Y2ckshdVTcS0Lu39jgeS1S8rpbd1p7Jwugw0gHcXgdAjyXo2N44RRTKWplFCwnE
lvoLxb3zv2llluhPACcDjsgSZf3tmEaEJase9jTJ2ldmuMKVOOtnaMSoc7rcFbGE7ttmofZzzsla
etVyHKUhYHrbmn3hME3nNxxEVP2e+GVwi1f7c+qtuPIyCTc8Smtnn0NLK3/B5H/LdQyhdSSTgQe2
+cLyZCbrekZZkSz9YfGGd+dPv+U7AJMRoZNh5ys7JYkCkuFsZv3vXMBvo5wEIWrYdHBwzpZ5WDwd
Mx1Wrs7LNG/BEqt+c+pm4vm53plQ94si4s8TEzsZDKUUPIYRCzNpD+RMIDaZ2wP3grz/flqute7C
dcNCJH9wjOJGNZq5IxYOjoPlHyjMGwl4TfO5NMv+pFxqDhsrDvTnq/ain95dCN4bdMUGPfFqC6GV
iGY+jbDrQFJJwFd7GAeIvc7vdS311Ch7PrViBAKhGYltfLpYqyINXYvpVnhBKJP8OAoCP9PhwZRR
7Dv7dGSGX0WCx/UnL/6lhqpiEyQE9NiQDzyTZ2/kYyUBqWEVmMw8QtQHaMmDz4UZTfSwqMKHvYR3
LIUkgOk0gnUJzso5TyLwn1ZMk57XqFOYtiAxFk4Jj6Nm9K7aMMXyecNJZ6rkAGSiCmRZLX2Ex0IX
2g5MfbroBJS46dc33tvxigB6lJuMzHtHoIBVb2moaPJqYM70f/K4Olw2sUXZmFUfScPxDeK2l9P3
TmiiMqcKK3/yQgLTmf3jsqH6uiai3Qtyl3zAG6pKCe9cQPGhbzZzNnut77kaJqJxJK6Hrjht/ffZ
C5muC6p93R49N/fGRN/V1UPBph50J9ygliu7pEmrDtmgCmQTHDmADTyu6lX/n+L8m+OYuKIwNDR5
DRlAYNr+8OhwopsYlIHDtFAXQSa2NccGOmkQZaW2Yqi79Sbqyrfye/yFq7OM0fnE1CwiWg9gKjs/
lTUkc41W4PXolIhXEd2wgZFsCaFMPh/fD3I0Mv4L0c6DzTI2AirrC3mTijFgKP/MLOirBJc8z+s6
JO/Dp7eGGpoo09EfDCVsVuX70JCexOw0wSvigy13dGTMAycUqFEqm5m2CnigRD4/Y2ovDcwXLQnG
VKpfGRSUi2W6u99j02OpnQ42ja+mqpYjjmhRqJH7HXKj1EwR9R14M2DwXMlvNuOtD0naliWAM6u4
vbqY9/JxP+IejY+N5CuAQHkdGKv0UZiSYgI3Yt1V9wcFSp7gMGZX6j4NsDesUu9CG1KKVVgT1CAg
2xzniZnZeZE2M+QqQlALTmSSxiT9BEn3CAxWbeoGRpqcX+udYMbGBVjr3hZSI4xCWiP3Jc/5v33H
gVXueSBbBTdAKHUT8f/1FMix7IN03U+yymhPBSKP6qE8j5uP5YJCw0VQIjbYhejc2DUQ91JRD9Mu
ef8ySrbaztxbYo40d9rBl8xWLqU9k8p+N7L5B00GxlL7rOu//KEJORaD7xfCa8vaGY2RmmMA28bz
/C2INgn8FYoQ2wYTl9kJPVZCBc1qnLvETLRBDSQKdTw91txOZb51EQBrzvCCCIMh7+PB9bZfyIXE
tQGHjw8dETzHsePwQACab5iX+lqUevAutbqVFszmBqnDlEUy0L2S5mIA8odY1EFskUDtZX0Z3a4h
uG0lbnF/YWN8PLnKjPBArZwNqXn6oADhfgmJj+DpROWTi/w7aOFyemTsvyZqwbxTSbJTA37NpHPk
gYcQAwdGNGgIBSp7hIVDFEV+PbSan3DLoLrDBgkyjR4tImloshof5KEko3hKct0q5GVX6lkWy8Xg
OH1qwCLZLKPqqQYeM90Qmm5kh2oCjb/ZgJ7RmdjIpV7Tw1/A/lmUNsiMt8+4ao4AHly4/oONXYC0
MHKws9wp1rLyJfC2FtMKdP+nWUiCtmAzLg92CQX/crjhBCvWhrV20TvEERJ20upDr+0Zpci0hzJG
j4dzcQF84n6ynd0IaSKl4JT1ByrSNjlBgIX9wpAMPrSOMBR5Y8+RkRVdKhQQHYYbI/1dEbgsDrpx
Ufe9Aq92J5LkwpuD8C9OFwnmROCTdlk1yzdyIhkX8bMyORJIYYZb7hMTlMzClQCy2VHyQnaqxBSh
ncS+g3mRftZJZy98j2/J4IxlvnqmLWWOOoN6zi5uz1jVx+xYAh4kA/iw+TbX4dGTyA3JugKos+2S
L0241Nw5uDpj5+dnbQcWwEzQ/4Ymd+5ZMLg08qA/MjuqmZkcNupjfiflNaYT9hYqO+0AbnQ82kA7
xQV+7Lq1mu+uPOreoLPfxLdLCD6nrLnVlaKhMMBaZUhLIIIY4yZW+5pkg3kUYqnvF6BkkQ65tnUe
WWOeSNtKxtvVYsqqB8K5TlhflsNvBlFCoZYe6ZbI58sL4wO+l32b5McfWeGiqha3iQJKMqRE938C
HTdA7180uRPKMvT8N6wGx7OvXwZ6R5FXoCbq+K5qI+ry6cOQCcOnyZQHgabtt2l0kChws3RtfK9/
6jhBKw34WcNrMB6j6T6FXUQ4FR6Gc15Sb0dRNpW5/YY9GNopS0XO5TFwmkxzIwFhhoW52KPQHQ9U
7zEe15hI4bsMmGQPAG7AlhZuhRS6JuYxBQqaDxoPA5VAycHq/+XV1PtUk/7tI4O+TTCWAxMquVBI
Zzi6srIY00NVchayVo94L3TqreQRyvllDgllVC9vGsGv6uBzmCBCP7+hkuZNRfQIXLx3Ym8Q94HW
Hg3ERPjGaz2iJmI5FwfmcE5ztehHMuAZLZCedUcEwdDXmMK3Y/xhQTGqwE325cKwMfvOeLoJvxRm
TCwLD8v1fBmnVjYRKuqpkPXL/0lJ/9/TKUO3af02HsyZ5pEctFHuoFoFS5GSYPlybam/bMZeIPj2
yqC4V2TkwFcD+CRXbed2f6FE3WbaTbQkBdOwnyRha9wkHXUpJoAZvIcd1jg8BJAr9ZZk3x8oabkC
ukyhVthIKpft+RvVky+TeujTzG089e0+wbLG50/+743/dM88W67vxiifFffH/qsohEF/p+pC5XUa
1T24XQQCIIJxwA5H69XoswdjYO7M+9upU9pHOwPXCF+tGDonq3vaRk4S4IebmI8fdMAmJAqtaqPL
p696dxJW2NFWYM/iVmhfEM8QLackUrLqkcTMC73qhU/J0AwhHBC7PFyDjA2CRcauLy/zr+tg6baU
K8AZKPg/oMakaw1y67vTeH9ESlPbVtI7dfGwPPXpF9dxHkUmd6gWZs+iPsJyPapOix+dN5xIFD0U
E1JAZ5lcl1+dHCEFDVPxdB865nejp0oHFabwgoT74tOJ9P+jgQNsg0OCk2VvZjAWnMBxcQLdyM2q
6AecGQTiOZCZEelpFa7dDYzPH81SSk0LkVVuXtVBJBY48GdEMXhCQ2GDxtj4Wpm4bX0+BitJMojg
7EENT1bnBt1eZd+t/rPqiW7rEplSXGQGtSAWAFy84T80bONWjsFn0wkCV4XIh+qDU6h1IphntmUu
Grm1MVPy6r2pRs96g4l/4mFlnYZwConP7y2ZbfHIoPn8Yb7t0dCIbKOx3iVcvM3IadxWG0MSYioN
GdeRIEjtNKKsddGI04DFre4KVjkhpuleVuxz151cs/q8/V2F2nDfwEdW9wciKlY72mPr6Mf52OYQ
UqBrOxMY0KfUcETHeirm81bWhgeCwd41KI9XWRon4Zfn88viui9oyCXRp7Ps0okyLH7XmF4nyRz9
KsNpunuX6/gzuIA26szSLJa/YSHALkA3xFzoyXKER5kLRBaPrRG2SOiPJKmR/qYJrtGZWFiKdbld
0mKmr0gDInv5UfVPEfIdaCliqigpKTRvElhU1cHRgPfpk92SouhwiTYEoyAxkIYmwbfe239cKauQ
ocS9CdSuOIvhxjxK8PNY+o9SaQb6Pb8DN4IRhfuqIcwfhp7uL8RX9M0V8gveJOYc/KSarNZOmun9
cu+gI0X+MfyVf4+2/7NbFNzrMQew23ncdwazsgKuAbWfAPRDMn/mdazlo3Q+eRR3XucrnuPXd5jg
Q/01Ouwp5qp6uFTt5VLR4p6mHQ43JcMbGta1APi3SEIZvG4rEJcjcBVD533C47ngYRmQdVaF9xzy
Ads6rwCwaQGASZo4RKbMhfMH0cnJoghbmaRN/hESdFAeN7ZxLzdgZmiaFiupKG3UtlTlc3HXJJCZ
vNK0dzCsR14TrjM/gwJIXvj04EfjCvlyvfK6RtClftneP8N3hg+l/hY0qxq5UAALjY3Yxe/h5+rk
zt0HXhhfGswg/X9ULjnOC95P4hoMHTuxxVVsCqsMMdO0jK8zA/AnUjkO3N4IFApjLwF+fdrYcNWY
riM74YA5zymFib2Tn5MeUnAmhAbOVtRSjdg2T8og1JYW/VsbEnfCAViHk/ErypA2FiBSKm6iFxwd
tfv34oQZzclzVBKg3VvdrhiWSgPEwp0SJZjNnVtffDC1vPIoW/ckzgbgOktCljXnA4Fz3qONCqAy
EyJvEgExX3/vUO4+QQJ5qM1c/x6KMgceQG5ZknAf5XqkEESDSwkc3VGrIcGPFFVCrdboMOyqP3C6
kbg7OPmZVkVlb7JvBJ4ksABdWO0sRlT4ZJ3Y9L3Tac9g6o23+DMlNUFOdhss7QA3/RdW6lKWAchF
vGXZaoZKAaNA+keD0eMZ9hQ9ir75yXiATtYcSg5i1xmYZq75hN/1FStyQ1heeeTfjH7Jv905V2Le
vbBjJfVI6QFusMJICRHIOjpUcHmkcip7ph9hHCEp6QDaWXnmYgU06RfD4SpEeiFKE+zfREHHPTQM
C+aYxc8mZBSE7hL7WducrWJ9mUBi3m83RHQp5U4Ezg9PFcO16tMwVtQdRWY9HeG+wKQwV61hwH8z
qTxbqJX2C6tdvu/6JU4e+bMGQ3RmGeKo+Ud3v9cfniUVBgdgd1F7FBocvo5WB10vVFCXGmFxO//1
CMLeKAQoVRYxjyeU2gkd+Gio3RBZhqWQXMBisnm2+DVfyt57QTIk4OYERfj9zVg9aLyqmYO5KAy2
mX0A4fPxVcDaZA2hALnqyqw7vSxrL9FfKOs6BNQ1B6VoEW98a69pLoaGOEqQa+zx5xlpolCBMt5p
gJjKWzJYD0EX9kaGtCNKQWrEPV8hWeytx9/EcGfWCTlqlVnjl5sdNdtv6jWZK8xo+Qpzz1HI71G1
MjOXnQIdKXrufymuuBzoO/UIdE1TkeZSg/gGWHWlDpWI2qlvjCxyPQu/ymdayjUR/yb5+Jfs+Is6
NTRg7K6KAKkyWgvpCsVdvBwL9QppTBB1a1m+m/EbTFnupsvkEC+QznCeLGbNBkVf6x0UDpJGWLKn
6Vf1EVQkY1wnbCVj8+palI60OkzvNjFNjHV7+1h7/0aByidPJdmDwimoBpbcMgTdMzrs01i3O6GH
edpxW33lPuLNkUh+On+nTv51R6q6b0oTUE713CGSgdk9wO5XJ9BwmksHGt0ZhXq1mV7srfd5n20O
eq8+NT15XbUhsIckTOtU1W6ItQNjJ6lgW7hOnWqbNH7OZbVED7ESkTRZheRYvyA99hYh5DJdHX9M
lqXED83cPMScwsJ/7MhSWzNf5ocr6f5ZDxhfoe9myq5PaefOxQRm89AeIQpQrhSMnWJ48ZI3fuwV
OH4uODYlgwuqsCaplKLuuB5pnAzc3jjfmSkwwOWVQmfSvLF4rEajvYw9nzOiJwHFPFKxWUC19W8n
Dt1t/W9G509h0NSYZIJp2L3TLxw6RgZn74JRoCHKMHtHER8RbvKrs8rtPPvH9Kd4r7Zo3IGO2iLx
Z7Tc7gUqb1Mt0b3W7mgZjRULUNL6d26DuHMLjDfKryrFrZBQF39Lajx7bMEnCIQn3+RukUM4lofL
pyh1pkY6XKHIsBYEEAEsPStSLaOGWjCsIHynS83nnhra7ydk5GW41DjjfSBmf5ErkPCyW8yw83Go
V1y4+E99+RMg3ccn16KW6/p+ORpmgtGsKScvYyy0BZiKyEJ+vytiZyQdkkBejw4qOFzsI1dF29zs
t1eHDyBkLgrwQH/Uz2GBff4sbHn78Oco/69CYoWjTVRTtQUTx9GFsB/22z7GdlJSulI6a0YJEO39
Sn8vUaZiUmPxHQXBXMmHzdIdjwqg6HQl+6OWgHaF4TdZaH1AGuYrdvyRYq4t9B6+xO+nQUBRkeoH
ZSJPw2AeGD3C6Rn1zvuj5hJdREitO8ldCHaiYRqEKE7nrzlW5RV2lckz26olmB+4p2gGK9t0f/TU
KIqjOacyvkYPAzx0EicIVVn2/zWQNfrkjPtmMWjXcVram4HVo9nn1mcy5n7HsT/gAt2GRs3IpJK1
z4CyEm9bsNLSYzlxQXy3ndT8SxxEvwBAculoAuM2cNwYNXe6dY4UTLlvkAbFwMMaS4o3tmtiMzPJ
MoHmNeHxvWmazw5pZ50Q7EvoukP3MU1zC0a5IGYcHniIiqmB/HBGcZgIjYPvX5GQMKEX8JeX9aN8
pehBIF0PhSx+Ok+OA0c1q2+DVp4c49OL4HX28YxXo6babWmjKqzOcbKUFnh6/YIKk1E3uN4NMhRP
8xO6F0bRryL6egmy+mdfiRw2H/Fsjk9uC49z7RVg9mNQl+M8A6J1ii52QiA85k2gkjnE1JcgKPJt
9Nl1Tr3Uhjr3e1lUyaZ34g9zvK+FYdHsDD/dnc3hapkXIts+bngrGh2ZfXarqDHtp1czYpB+CIXj
oT4mGqvhrDIN1rNbaB7LJEfN6G00muEEa7PSaXhJ/SwBL0tcYsuLLF4iTa9BmuVu1jLZMy0ztQ26
RXlr6zwy9LGS4m2ryb2dK8xia23WBgPJ4cPOYiIm3qD0/zsZMWWCiIlKl8j6aH3uXk2p25/mMipX
86yGbPyv6Rd9eqlTVsZnnOFMhVnjDOps9p2KVMvaWQ8TXXmJz6N0rS1YY2nf00s0m3TAsCXRTmBr
UJxkEA3pDNVTJ1d8JLCBsb6WGWDbWPd0UR6NFM07Vs0mRRxaRzu7seRtjalxV3Nj3WQO/Gsz4upu
8ln6FpqrAmizFZDwurcH6HLlg0r4eAeCfguiHsVBsmsHadxutcHlWIdZZrbGIzAsdh0cbJ9tFVOe
UTDMMB90b7oLWxLGvNgc9AyuRdHGRYyb9I8OLz5nPN+46RRUUR9BZEX72KNO6EH0U48ZwDIfGZO7
0fBBgKKUumVL46MrHwLGVkW4WW+rfcMSYJs3WamCmnnIltqTYctvS0Kq+XngcMiqOlPFrJBs72hg
DwpyliV09Mddq6+XdFUiiePQmfmY3mridpWscCeuNkqcFVVcizXNbhMq7X1NjdjEjlcDB40j75MB
bT4eq2GaI0qG0U9cWOiAtPmkxs883nBw1S0SJ023ggEXVsHiVKld9zE0zb8mQYXBMW0C2Ef1RryF
bQkdZ3BKMuHLBWzZ8CGm49j7uxcwjshjELe21MGOkTStRabNi2KzMH6EgkE7wM6eNHzreb1XD2A0
GXREtTc86RQVRp4DgSkXmYth+1J5gIYkbIrh9LD3lV2WoRsdpzAJiL6abgZOAu0=
`protect end_protected
