��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7�r"�㤞��dY����D����0���r[��)�iѾ^�>3@hI�2����kװもƒ (&z~ͦ �IU|�C����0\>�\J�8�UoO�ұ���Tg ȕ_���ȡ>e*�/�}eTE��d~��n�\�h�+og����˳�,6;�8[��z@�Q��4צ'�]�`=Й�˛�6�Ø���O��BG��4sU�e����Mq=��w�k�����h9�o�u�U�qD�XtՉi􂐁r��H��_��wW�����L�.J?8��64�n����qt��8��� �]�%oh�}iZ����M���M�1dXnP���b�Q�K��ض1���M+Wf0��˔��P�E� ��L��M��R�-���rkj�^�{��!�3���f�z�$�݉�Q���j�X2#xӱ���M�	�"�c����8�y�~9a��}]�7W~�F��O��GԾ;��trM�� �v���H��S1��-���{�}{d7Ҿ�w!�fc5ύ�(�0y�z09WU�b��QH���Y���7�y�ů'r̩`���������g�:�V�?���F�/�^��·�K�<7 �Qnxf9o�2̣ef	�fcfr��T΄;zDY��cNAE8�1��'N KX��چ�<B��M���RS���ݦ��	<������;�u ��k�9�_{^�<��V�@�z�a����?�Z}5ޝ�nx|��D�\99GQ�w�aǩ��[��p�.?e�߸��ٸ�Q�p$j�a��%ޘ���&A�j��_�1nVkƘ����n���� 28]<��kȣ�U���䅸ѣ_2
�<ВkbD�����{հ	�� �+´��uw�H���dn���c����S�e�%��ED�3�����Ö��C�v<����f��bC4y]Q����6�?���a���i�H�����e>���/���A�6O�`,7�z��ׄ�������m��pa;�!�K~�,�2Z�I]���9�d��`O��:e9tt` E����=���$�k,O�M�ƠE�rCo�9���q����U��S����8]�v��bw��$��"[�08lߪS�-��)UC�l��N�r	D��Z��)6u������V�D]�����d��W�,��&�b�y�f�2�1�m�7���"i�z�4����<����6��1K��T������5��F��!֪*���U��/����R5���jc�<y	�VD��|�3�
��ٿ��^fɘ/{ �:���=�ӋJ�*
8ϱ�p(6�|��۱����;N\�9-(�D�kMkF��G��� �bI�������s�&ux�]%�Q�`��w��Ӄ�Юt�Rǹ�$5�=�!���&�2��g���l�xg"�@���c}�����rO�!z��E	!��Vݥ���4NL��ruRt�JC����t��у����O��2'S/�/o0�����]Z�:��~�H�%K[`�3 ~�e����Eup����BP���n,&�b����cU4
F�CA$W�!���$VG��%�B��Y�w[;��a���������L�(W��A��ﺧ9"
��m��; a뤫g���^����X�c�r���8�zxa�����6�)�/�Q�a3ʮ�2H���s$���ҔmJ����8��W������KLq�x�l^1�Y�P�mQ�}$�d�%8�f��R��@~oxW����L�Ө=�$$�3g����e�?��]|��(����ś�����!6��R�uWX�!M�]Z��R>_]�� 7��g��X})6ZtU��9�p�t��s���0���A[���_��3A͝ ��3 �-!v'vڏBa��=��=K=v��w?�9r"�&[��D'��0�&��W8Ԕ���LYʆ�wl��';�������X�.�Z�THK,�#!s�� s�}P}���ف~m_9����������I�<5;�E����}�v�$�g���Wi��&�)�4!�Q綟%J�)�i��.]����u����i�՗�~7j{�X��N��q_u�&��ۈۺ�{P-~_~����Ƽ�� =g/�d�����wmJ{z]P�=���y�Q+��봫.�F�<8L�!A��T�u��8��k�0�_z�����n�fm1�cn�t -�H�ϴen�8�B���&��ȰtH��$qH���\ܯW�{-�CI�����	Z�9Ħ���|r��!�j+<�\8�����^햞��E/����wHc�]姴�B��e��c����0�g�,J�#B2"�[���C�݅���ݚ�u����D��}2���-:�4���R�!��[�ݙJ���7,ʷK>F� ���$�)��������):������#�y��ǭ..`���<.m��߮��� u���i��b��#7qvmL	** �Уf�#J�!S5�� ��P�	�'�6�ƂN�7��*�"J�����\�\j�~���r)�,�ytb�^��G(�i}�^TJ �s��K]e�z�+��lӉ�R��$�}7���@�q�#����Xr�˝��XI�W۷�d��Dv�C�ih�*�ky����	�Ҥ�Ͷ��L�'�����Ow;0k�E���jV{0ڗ�`���W�D�G_��~U�_zԧ�}���W���COm�_�H��+"�K���?N��:ٙF��N�8�j3{�uW9H�"����5&>�P�_�$�Bb��?X9�a��G�ȵ�&َ��hi>JE4��V������K��)1ס��%R�?y�1�w]/-��J���QU�|hb9��L#�r�%'>�v�Ѽ��O��L����������^�I|�)�G����	�.��Cġ�Ҟ����T�l|3V�!J��#�gF���?	�����㋃���"�9�s��P������E3�Lhݽ��Q#J�n��P�A������8a�g�B�&"S �r�!�1~4y$�د�4�4R0#��v��4���f�6��׽�����*��{T��;�G��b�Ѹ`�+��1piR�/���=�*)�?�R��~��(�1�|0Ӥ� )A�X@��Bt��m����gn���UW�K���8�@'��^����ࣀ��������t6�gFHZ��{�2�f�9�zm��Cx�����1�����{	�1d��=F��OI��O��ʣw�ϳ��Gnl��	���u��w)�7�b�������}�Ի[��?�J�ޢ�Oc$dcs�Hb0,5�~&��fP>�����â"��7v�1t��+m��)��>�\?S��-�Z$�G����qr�U�";w��%{��N �y�"���-9�;�5�<��V6�ȼ[x;J��?7�&V�@�怴۲��yga@������;���10�
����Q�4f,9���;V>�ML
HQ�:.a��~j8s�Y��]����!MF�P�`��}��8ɎO���.i��Ο���_=��A��1���T�Jh��9�?�8
��ּ�����܆ge��-tҵ݅�I_��H��i;��� HEw%v�hIC��F#9Ê0JW�[x���Z��Ec%����LǨ�
fB����B����*1˸w6����O�!3��#�E�?�>�f���q�؞!X����S�r]m�NP�Z�k�?b���A*�香�CSS�J
ux��Z��.�U�Ե-�yR�fv��b�ٌѼ�~KKU�^���`���<�q��$4��[W�Aa�u|��(��-�{"�T�D �����Ŧ���V�M'PbY�n�\0L�+rheD��ZvuJ�;v�Jib(Eɸ���>�<%LqKl��\��{�_��:�M �|e��{�nv�I�$� �1k$i���q�Z����3��{�3Y�Ès�Ï�-6�M�6�A"#j��ˬ��"	K)�W������,�!�(�}<���d_'�g�^���5�ZƟ����g�
��8�B��>�>Ai�I���=��q��ƿ��Ҏ��O	�����s��lI�0��3̻�iHꙨ8�tf[�snw�������ZJ��
Gb����cT)�,�1s�I���c_�#;�\B4J)6��N�̊!�{�R|4/�To-�_	�|ܛv�8>dۮt�3��f��k�I�j�� q��[IQ{�s���dW�F�4�������V��#� ��	@�X��F-b)T����3�9{;��r`?�k�-���K� ��#�4:��,|�K���q��m)���B@��觤:���w7�_�}��Z����.�N?���V��(�~�������}�\-�!XI�PJxTo7�������\A9=�4�4��ʖT`\g��,�79�$�:M��։$�:x��o��,q�O�QZN�]EK�6�T?�ەVTu�C�r�e��p������͛,����kIO�p�W��]���j-�i�B�Y��g_Ś��xF��Ƃ��?3+0p	Ʒҋ�5*p�Y�z��I�4j�P�����Do�����QIhȺ�v���>� C�V0����D��_�&ˊ�XD/V5�zD���bk2b�����Q��P�(�E�DFٍ�xBY�H5�O���لV���j��0c�hx�a�Z�T�£-�\`=��Ē��͏�V��Ie��ە''��U�k[!���ҊF�4h���U���N�0�NB���BI2���>3�)�s��M}E糗���hT�� ��M��)� �=�1�6�pZ�����؞���
�ׁ�ܾM� �s�á1��C Q���c"6�w5�=N°�5�F�n�gL�ݼ\G=0FpE��t���9�y�����^�]�� ^<Y��eG��UߴӨRl��Y^�a��ȱ/���O�ʧBRi�1Y�� ����v�nk�.u0	(�}�~9��8:��� 䣗*XZLZ|�1�,�D�"���/��)5�m�NQ(}T���V�n�u�y4���o�<���{w#~h7k��/k���o�_[��3��U�H��I�xk��{sI]���ޙ��>2|[̨r 4X�
��3�A:��R��ܳ��O�<M���=X��X��3�]������@O�Z.D8o��.>�O"Wq����l��V�}�8,�묑�X���Y~G?������D}q���W̾�>�ݱ���E��!�$��!��{c�����~f�w?�cA��"l���#A��gQ0o0(Y���7d�E	K���-��#�>v�@'�O�n�Gɟ�������Zp{YC!J��V!�NyI&ik0\�J�ԑ�"���3O����7�jn�Qs��S�o��i�
�]�����S|�˼R� ��`����5lϛr�N.�z����JurcF�Ʊ���d��p���4����<�ē٘KK���*�;��=�M��E�3Y�$F+��:U��B����u�-�:���>�a�s�-4���X�֥��dȏ����#Q�p�'ˌ0�9��.��xC�i�����0�b�`0�ߐ+��a�4��z��H�H�ٳ�ʓ��Il����w����*hF�g��]��*�+��l��&s���מ�US��|d�r�?���]�k�]4�[��m��>E�,)�ă�H�â,?mq�k�ۣ�$���A�w�C8��o ��ða��.�v�l��-������|���Ŗ�L��_�Ҋ�]۲��! �;�Q�������r}�T�E4�������:Tl4�"E��ǻS�[\8�	��o���RN��o����|��d���j <���8|2�Uɤ9������tJo��$�S��f�[�}./�,�l�9������AQĮ�Ҁ�iXY'���Č�������+��i���]l�������& A4�\Wȕ%MBM@��^M<�}�81uj���$��݂�i\�� �hu�v���Hir�pf~��-Q�L�b�8�ɂ�ͧ�6I�b>����bk{&�˛�ð��ʅ�j�_9r���{"�<����#��:��q�F,���m{/����~8��^�9�PRe��#cč�j�6�0Pvr]W��`E��i;��+Ϻ�k)l����-4���I/Tbh,\ʃDTw�^�1�T(8�@k�u��_��}��Σq���.�EݤrfB�7p�O#F�m,��K��I܈	 b%�jK�g"�	j;��7-�S��גŏ�&�u�D�41���#T�f������p^�b[>����@����6�1Dc�D�A���Yږ�"\H�b��h]�\/�6������z�V�)���,���<+�mM�zQ5�.w㹵���ǂ�!1�Z�:���/z8WW����p�^ Ex9��F��r3�X%>��("3��&��EIw����D�ke�]�w�S}%ͳ�
M4�|�E$sN�C�%��Psܽ��r!F6���|Q���X4%/���Y.nƷ�R�I;n�y�pF����1�$*�,���)�"}��T[7Sv Y
J��ÿ���D��>��{�$;��҄-�P{IK���B.+j��aK4�����wm�V�9Ew�Qo1o`���Q�<Y�����-�3[,c[�K
��isؤ�����k�ؠ��U�i��?�.nҙ��*ĩ�w�R�.N2 ��6�IS��F���N��9J/a�>�;�U\�8$�HXX�\/G^�\-ctvD�����貯�iy��@z��z�܍L�6Ї/&�S]L��dq`�11�CBM~�y>���@혼��?�4��ή2�{ ��М�6WL���1D7��#���-���})^a���z;3ݮ������;��>'�������!��Njv��0)�^Anؙ)p-`{;�q���b�/$f���3-KIӁS��7��uq~Du]�$C��K��ծ>�,y�p_�sw����	�{���a^B����1����9��j1sI�q�ϥ���o��$)�&��f�C.�N��y�{E����jƇ�E�+��<ڬ�M�ن����
g3��s��y�K�8����RU�6g�-��j�In7��~�~���ҊiDͶ�^Hgql<��x}�|0�3���X�o��_h�$�Y`D((Z0�b�?$�P�l