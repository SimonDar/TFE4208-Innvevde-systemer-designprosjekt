��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U�}{���ږh���z���v\��X=��΂p�Oc���s�?�q\~�>��o�-h����^M�p�q���t f��a����~���@kĻ�t�t��7�s�]�@G����0�땆&'p�T���s�h�$.���B���qpL甯_ʀ_��6�.��%��YuX-6~� %��"����ZC��ko���[�)clOK<��62���������?����ߏ@E�+
��=SU3�M$��lǆo�
���2��%�'�zZnWH���C�	gV��K���Q�����j�������W��0��h;S-��|r�d*��ּ��R�ZB/����6��R���?i��q�A����/�afi��l�?�Sܟ%��Y����-��הbm�_��;Q�qoa��}��Dg�ScUC�~��()�q{?r뺫�H�XuW$$�$��%�`k�'Fb~�F��;C>�-���02�ZnT�-�^�ﻱ���(�M�:��Fvt��Q��\��Z`�����b��+�B��V2����}�u	+ZT�3Rf�)�}�D�,��ʼ��YrEN&tۉ|�Þ��|d̥�k�7�j�r���C��۬�����R�[����V��:?LQ�D�b�#��6ܯ�K�˽P�֬({�RsO�o2h8J�������}�z��R���	������F�`��Tw1���C"�PCm�ݯ6�|�J�9��z.z��&�����5m�����>�TSC�����CkmErGY=�S�_S =줨�<��T���w�I������g�����`�Uk؞�rWU_�9`��aj�i�؍�U�UT4z1���p��y�R�#V�}�L���w�]�1%�����Z�-gy�C�㽨�l�e�pr
Q	��:A.T�ߕ�T�/�ټ<*C`��œ׏�Ķ/�W,��ӷ��B̲`O�Ha���Ҙ�D��֖��jl���1��i>�7�(ռ�%E!m�z8A	1$�'p�A�
�2��+n�h�_��csV9:���n��vGkx���N�L�~!�#��-���C��3�鬡��VKҌ_*�ݣ;�{E:��IYQ���g �C[��P������f�*�e[�q2�}�4 ��%n�&8h��f���My����b���w'3�j������@�~��\�s��*�XЧ���O��u>�f.�`��B����V�ʅA�g��eoZ!խ�=�� w�l�ߡ��z	�6�Y��G=�g�i�t��7����+E�V~��Ԧ�u��=����c�s?��]r�b�c�u�/���!۝؇[�P�*���o�h�؛�b)l�z��V�n����	��,I:[eo$��`���~S��A��H���|�m�>�ߝ���$(���w	QGB�a#bW�d��	�072be�w�~���I�"b�=��}d�wR>nE��A�c+�9]ӼbĠn�� L�}�o�#�sL�MY��T"7׹̄�H�f��8sTM�K��_�8B�r9�� �LY��j7a��Z�*��1��,��
~��=c+�͈�SC�5�����#���'߫d���/�C0�Z��qV�������9앣��򟤋\n���Z�t�K�4�4������)�e����Q��j�D�gm��LJ���ӖK]lmL����u��;m�妘�	ؗ�v��֕tTG��"�/��N�I;=�����R�� 7�Th�u�6��I_�b�gť5��1Ad���zb)4�o��v�Q!c\���}4{�
 �:��d�9&D?<p��ʶ!��D�^�����$q��*�v��>/�VL���~��(��5l�d�V7?cQ�o�	��o.U��Y ��B��s��
_�nQ�IN�̖'����<�r����U��y��S� ��5#v(c`��Hd7>�f������x����m�+�����&�P
IBP���Ӫ_[W:����.h#7��6��(m�!<�hA[G��n2���hyb������a�6��u_�'}��n�rX���X��Em���>���H��*��^��n������k��h��ky2}�1�Н�k�A�H�n,3��K�2�J�D5�.x�˥d�Ͽu�Kᾐ9�2Cρ�� q��!˦CF%k:�F8�����^M����$}z� �{���-�+�A�IN��;�Ლ�eTS��>��O����o��2w՗k{׵�������X�bG��p����($�^ؿ�/ĊN����({8��,�$�G*T�[ �q2��	���Ъ.NrqU�s��������b���
ȯ�ɨ�J~��qW#�)��0�{���:H_(�k��9m� 'K"	����k��ӳ����Mz�2��a�Z*K�:)AZdy5�K��2���;��/���v��r�Q'P�s4qԎ:1?q\�_Vw)�?�=��
����X�s�4o{�GR��w�⮍A��+��.
���QH�R.������訋��9�;��؈���WP,v���Nŷ�O g�ɨ1����;�n�E�W_�~,4i�bC �a��ZHA ��M[֗��4�`�,��/����0K�W��p~���XGP/?PJ%{���Y;���t��j�:@`ǭ����!aL�! 8D�"{�����}�<i$1�U���?�
D6}Vj��>'��&_s��'߲���l�
�qM�=�O���;�ޕ�^nGk-�y�`�N��U��m�I��<Q٭
���x�X`'�w�$���zV�dN�c�M�V��?��jh;�9o�����S��	w}�fiP�.#�&5��1a�j�~�ϕG��	5�6�I���.���p�?D��,� 4�:���p�F��Y�mq�ﾱ�$��I�$��c(��Y_,xz��l5�1���.�f�fx�eh�/���F�������w�zz$� �0w��e�Wi�m ˹I7�UM�K���+��<�&�!�~��S,���H��B�7�v�9�TV2 4�@
���I��	�$җٺ�pLÌ)��NzzR�&�~P��]\։�˂ȪJ�{�Q��ymj�������V�u��<�n��A�����ı��$�x�6��l6.7��=Nz�9�..x|��Q}��#���F�tWxäS�=ۮA�n���-�r����]�K����0}w��e�p["P.��9��vLQ�`}/��O�����l���$t��u@kșW�E�*	��y��A�v��q�Z����[m_��&�҄�I��'Op�I�����M��L^A�{���ǯ�hc#I��q�☼�To��(F5^����9�a���l�m�|Wk�_�R�: �~�^���������O�X����xՎ'�6�\�nc[۵<M!@�^��穢�c%�pb�_gQ���V���]�Gm�a҃xn����?5�P�뫓��)wN��l�.�:��i��6�(������aݷ��m������Gݠ��4W��vO���i������yS[��X�e͹:�Մ�i�K�d�i����sj6�s0��<.�4jfK�.�m�@9BZB�Ue�b4�j���>Hy���
���
�IN�pgcmO���g����:�7^�I88��ވ&��`��J_�����c{ӂ#i�@/�<�u�B$]E�/t�|����H�L�^�~�|9�Ԡm�k�(�`�j$Fzٟ����"G��;����M{�q��@683���[����B֝^J��)�E�E��6��F5Z��#�M�B��
�(M/��sۇ!~��l�x���]f�����x�,��W�IWutX���}O]��L3��M^�h��
��j8Ü/�0h��(a��Y�x{��.�
���Hic� ��1�]���ء�8R�-��s���d��G�
ӓ��-��ڤv���?�y��L��!ir�	��-rz���Һì���0d�s�T
��J�R�/ �� $�5��{:Q�G0�vWA�C)fJ����efE�l�>�r{���>H�������|�0�R�$�������Q�x4}UM2�D��{I)��S�Z9;{��UK�1j�ik0;��g%�S�b��L�ǩ��a +�!�n�%٭�`�%�$	�\����nmI�p��`�uF�����^* �@Z�<�+�mf������ܢ.�_�p��j!V�=)���M�3�_�P���gxEi^')��dq�G�IF�}�	,O��g�YT}d�Ɵ��u��P�!��lq�:����>Ct�z�À�A�A��X��[�j�s�����i{J�(�-ϧ�ܘ_	�Vm&dx�������i�^�-Xj*T�Q$^X�s�t��mF��uv��j�*\��]	\�W C���0��$odO��Ҩ=^������$>�խ#��Ugy�Z��}�M�)��|w��XVt���̘Hj�/@sjv�!�ϥ��m��f�x�^�Ì���M�V�:�K���2�
x
e�vg��;�Fm��L�w>�⓻�����#���ə}a{I}=|[����&h.����_�п��U�8�X�H&�pz,~�|� E�>�49��&����o�c����+����p���]Bt��؃�S���D)�����{w��)	|N�JJ7���*c6�5A��h�
F^�Z���z�:�e�IBⲆ �{�7J�fr}[�
Ú�)loܥ
�Yx�1�߈��\dJ��+$�/�y�{ �1��&��i%����� ,��.�'�h1���(P݃����ȴQ�A�U�+��ج&$/�Fl�D���L�L�W~ x�j*�9���hwt�*�3��al%ѵ�jQ�|<��W��ԯ��)ˡ��'���~,��\c�d���R!ӹ��$.�f��=v�T6uJ��a5ܱ���Cq��A<I��j��xL5s�N��kGJeZo��ݬ㥧�k��avh��h� N4�A�9�C�J6U�)}���kqN�gJ1��		:� �͞u�6�) 	�ʃ�z��L:@��6'?�[<�����g��i>�_|>ǥSJ�ML4o���P-{��w9�Qy���eW�&X.��v��qZo��k���v\��|�<�P
����%�E�Y��H{!�������Da/��7�B�j�G!�0���ͩu$�g�mL�=b�����p�c"�[c���Fۥ��juU��W��R��8TX�>j�8���%,)`C�$c�K�t���
(�����|�U���N���� �y��[DE@/��a8T�nA3� Wt����
FE@af�h��ފ�)S�[���f�|�%&r����.	��s?͵�Դ\Yr"	ne�qR!^��5��	ڸ�6�E�C7Մ�,
��up��Z�����|[X�S4W�8U!�)f�y��*Ҏ�J��Zv2�Gp~p��o;d��ɯ�d�]���U�^l��J�L(ؕ��L�x��}ۋ`-�ҜE��yX)��]5/�e�Vܭ6|�֠2��`��?��Յ�2>)9����@�"�O
P��*o���Я���r�-��E���er��(f�>�@�#a����L9G<��K}��"H�� ��nc'�S�R��N6 e]��z��}��W�f���S,��W!��߂*G����g�Y�3])�8��rw�g�n��Zgj��6���=�O����Z�e�Z��6��oM	a�UEoh/���5v!fnԴy����y�?*�6ݰ�ϓ��/:��Rz��2Ԃ�L���{:K�"ˬ�`}�@����ܢ��L�jĚ�9�K�	���Xk��Yo�K`nG>5��\M����"oY�2�r�6� p�m�
=δf������~'��Z���E@xئ��i���<P,yG�p���I�=���\غ)>��]������'U&&*��鋮Oc�ݬ>6I��v��G�F�!Eޝ����9���$���9��7�{3��n:��ְt��F5jU��ZX3��	@�Y��U�D��3w3?�P�_j���p�ͪ��O�Wr��&e���T�6}s�
w�e��}~��Z�l�1F#8����\�}�&��*�&�D�Hy�<�5%@�y�A�(��&U8�q�L�r����V�HB��� Ã�3�β��u2^��`��qƏ��ҁl��dw��X�t�@ʌ�g��,s��X��'lZ�j��1:�_�.Bpε���ozW8�5���3��r�m��	.�����ݟ��}�c{�q3�"�%�*�D�O��N{�X�`�J?)6��)�x�JT#O�Zݵ�i�6f���b�G2\YH��n!�2��~�k�)���T`�q�g��U�"��T@����gn�]*oo�5i�xpMw*�l��@�Xw[/����`e���	9�vfZ�Fﰯ�E��N��Dݭ�?�n�ʚ{�no�\�[.�h�ڶ�a��l����Q�y�ts�y[n�1��.�q@��א�/H���f@�0r?3Q](x�7�cq�z���.���������Wq���1hs9�������דs]��T��T��if�1�~5%%����o�$��Rykg��#�"�	A�8&���2��g��~b[�����M��q�ˤ��zx�5^WG��!O�}|&T��p�B�6M�o����q���2EY^�c�HoW�$O�U	m�7��1H��v:su�� ����=�#����wk�oo_��j�#e�z��	�����uӬ��Xp�v~�Jm��'����'�T���`�  K窃�<q[�кDK/gd�Yjc.�������\/b�3,��]�z�2ڙ��T�!��N�P):�����(�Y�R������V���s�5��+d��=���I��2��8n�H�T,�D��9ۿ�Z�����b'�ǟ
c����J�1�����(�#~�,��W)[���G���E_���gਖ਼��E�u�y�r�}I��"�|�݆���5��_n�d���v�p��ULz� Om�"��a�HX����k{�a��FM�G�n�Cw���B7/�O�j���nJf�P��������+l�Gv|t1<"Ұ���Ȱ @[� �ͶrPdj�!��}s0/x�h�y�;z��gµc��|S��s�*��a$yt.:U^����gl.VqC�[>����.zs�La�̹b.���Tgã�����?��)�k�kǢ���7l��2qDTMHyY�"�WK��H�A��Df��<2�&�&�-�D��0�n����Ax����W8�������菠|0�	�N2Ǵ#�,k���X����	�/�0_	�P��x�XΛ����jX���u[�'������ŀ��b8�\I �[��R�D.�gM��KeN�1U=����Ek�S��8��R./�>����oL�ɆD^�r>b��0eGJ�+İ �B�*�B�N<��X?�q~�ce=�"&��r�GoD��7�1����:�[v|��v�G��� �2Gχ����4'���d<���WX v�I�������&2���� �tC�u�,��'C}6��p���&nnL� c$��b�J(�Gz�W�A�j�п�����0��S,��"�܂�����s_w�.}�h%�����>�bɷ���FE�f}��cH_#�����`	����%��7^�����P ��f�&���`�|z����p1vy�s�?��
L���Bh���̐gRLl�a-���"q�Ea�X���l)7qz���@�ͼA����8��R����W�ؓ�#i�ӯ��!�3����B=�!4�����\�����Qr���2�����u�-bk�p�FL��GF[@9}�c�A>��'�������~�lT���W�,8�7]V��"��]�+`�;� �bI�%	��������x���G���WQ�z0&��m�z��6Ġ%���S#��c	�������cZ�z���vBwm;%)��(k�A���sJ�g6�
 ��sd>���<or���g���z�z�� -�dCb;zɕ�wH��Z6Ў%��w���u9��l���j<93�MH{@���]�me���lj��h,�4���Ja��K�fp�� �����l�����0�e����7� �	P���o(N�*���յ����?*8�[#�b�4��L&�ް�͕�ss��jU�jB��R8QViG3��~���#p���j��J�9`��bj�@����8ysR�Io�4�M�ݧ�LQ��&`��z;Ĉ/��;H�W^M�J�,�_ր����q�e������y!��e��rv��ٴh��Ij[��I�MΫ����[��Ⱥ���ש�	o���k}�	�{��ƞ�T�]a���
����Dͼql�6u�5�+��5-k舚yQ!��1�<��MNߺ��IaQ>�51�����J��tL���
 UX	 H-XnZMg���|��[�Q ��΢�q/^�a-�9�Pj����^t�O�����A�Ju�zY�9#Ae�&��������Zdڏ!����
Y�̫�dt� ܞ�;�2�v��e�c �.�_��jB�r�6Ύ�:� ���P�)�I_G�֞����80+��$���#q*��ms��2���+#晴�TB ���0Bd+m��],�ҚK�-��d-�_��78���8����
� ���L��\�<M���	
����6I!��]�I�?7��6Q�|^gsJ��z�/Y�z��D�;�"��Y��]��q����A�;��8����AXP��A�{釁�఍�ԩ�g�a�q=K�ٗ�\���w�������%�r��QL�4ެ���<��a	CE���*~`��Ed��>Xܖ�^X`162x�4���i�6�Y�k �6b�H^�-Φ&��^{ MEȓ4ˢ�m�� bM�b_<���7��PW2=�E{P�	,f([	��컅�-�9Q�?���*"�?��)`��h/F+@�¿V�Y���_Z ?#@g�2�tǣ���f/Bfm퍃�7Ts&|}y���᳙�e2*C4A�M�0ͻ��(7��X�I��m=���\�nLp�j��N��[w�6r�Y�(�Di��R�J.��ϐX�>E0?[��<�����j�B��pg������T�˩���h%�P;Sh���~�Y�{��e�<لQ����t�f���@B�&�U��D/{?V�-,��Q��*x&�y|x8�ֆ	��_�0�4�Rx`1.���.�C�\d�0��i�65���Y���a�V5<{�i��X�w%�΀ �2��]s��(��(՝��|'���"�q <�5�F�� ��lRj��
+CK�#�u�+b��a�RpDa�:>r��V���a�3E�92���f�����V������	��0iaC���e��=�j[x���ij��Z�xm�4��'t,�`ޙu ��ϧ�M7�
�� ;���u>�=9�"`��HT��w5iΖx�<�(H�#��Ȟ���B썔@��Ȫ�*u��KU��?�<����Lq[��o�#?K��A�x@i�nܑ�_�ڝ�nui4޶�:��5��	��ھ� �"�>�õM�n�P��� ��B�U���#��<�S&8�X�q�Vh6���ƈ��0W�T�$�o����c��B� ZvF�[�Ϡ�D�d�7��2� '��LD�0����R�i �C���b信���}2=�`���"�a©����+�&�����FyW���d�0��!{!nw�1�2�X ߅�5�*[&�WTM8�+���<��C,d��t�� ��Ⱦ�	G2�e���g�iV:K�䐡�}#�'&��m2&T�ϼf�FR�U�M� Q�IϿnļ���{a]v�F��s-�ə��.���p�fv4>��s���!���q�v����a�2dڣ.�s�����|�����{�gn�a;Sڑ6��J�����\�!�3��|���zi}sC��Ϯ�~��y��|i���a��2���/����U�'��b;��SK�S��'ғ��59Y�~�QV���@�l
����[��5�x��u+�5��=��z4��#r�I�'c^D�d̀�c�j�B4��p�M	�[ID��SW�J|.X�m<e����-T�vV.��\]e=	�],�ތ�?3��� 0Z_�+�77�ҳ�"��D*�dE��/r��h��c{�k*O/�?�����(3u��}n5��;��g���O\BI7AIY��NNlH~�[�y	7����x~}A0c	SR]��~t�����N(ּ�㑜��(e�C��~ZW��O��Hk����� �ds��s�"���t�������Rl	s\Dfm
�k�Ds5#��J�� �Ua��1�~�)�mL2d���%͹��W�4nD{]x�@+1�t�E|jk{����_��B7I$��w�0�YO�Q'��� ���z��Vd���X+g�xq�Md��-����K��E�^.�Vm�R���/�_-׷8	BX��a���ԅ�P��S6����?ٲ��Wq�!��r��]�"T��	շ�)F�!��?�<@�9w$�ہ�ڋE[��M��7��H�1�t���>�U�W��uò�b�z�A|���o!GSw����0�=c~wi�f2Α��N2�R��!�c��{� Qr?-^�ѡ×ǁyr����a�&�aq
c0WZ�b�MsR��n�> ��Q3�G����o��D�����H[��E�/Y0t��l��y�D�%�{D�o���U	�o˝�#�8��&��Ӆ���t{���*�lU�Z[��^'�\kp�fA&K0w%����2}2v���E$0�����I/���ǡef��v��5�!]3���رD��<wg��L�@����T0A�`v�i�\U0�dc	eOvCx�Ի��m�OHxl���"�@���僱]����hS�-� �=26�$�<*���5�G�h6p&��hܰ�p���Fv`@��?��q����@a�z��+*Q�;�vQfFԁ �dy��e�	;��{9e�v��il�A�~
��s�Zs��,��l��M:4U�|媠���ViI�:qn�U���刦fa��Zx#珺u��ށ|:䞬{r��w����~�����V�bKK%�k�V�i�TT�k%����]#���NH�z��
�Z0�D�b��_i̸f�KX ��6��դ�{�@|K6�Z_h��;ln�8Ċ�i�n�E���9-6e5����[�@S_�Ą����ٿ5�fa�����vkr@'d�`��c&}�6k6���"��'��U���X3<5��?� ��5����5$IB���?q"~��DBu� ���sB>G�ݿƖ�(�J�#��H�h�̴*��{�L��F���=��恽��f�:��R7��*�R�ma���a%�;��̓$U���Z.�A;����XZ�܈`X����y�����8x��9'��z{kk��u0M�����1�}��w\��f��;������Ѓ�����"Y�iaF���鯽�Ú���t�l�Lu��^���s� ���������|�QD�����`
��3R@�� s���{e!n��gB�SĬ�e('�J+�:~fF���=�p�`M`�h|�6�&���ٟ<���9����c��	kڛn�7�����s�`�U���-Ն�xlhb�m�M�P�^(��\2�/&Ƚ;2 ������AQ���(����y�.�
[lv	P؁L8����4l%0!� �<�¬�m�T�nZ-���	?�g�D���9N��u�u��X6���M�����S=F�7���?a��A�`�
�����e~<��݃���·�ܛ1�ZvI��n��ͷ�����;J/�T
��	���
���i��)��7�:#>_V�c?l@�|�ɰM��=)�"%���G��5�(�m�f'�9!{��2���O��0t׷6��[K"B���7����m�ﲳ�я���UC�x:o�E���錐�%��a�6+�T���ܨ?H����}
�.m�p�uWup�M�ԮO�@�O�@?�����FV��R 4�ys�E����@lPQ�����*踝�IQ���D��+� a�Z<],!p� �QzݙW-�.V��Ż]ĝ�d枴�E�ēj��VP:�����0�`�O0��$�o��zw,��o��I�k*�z��a�n��f�0��Zh!�Ղ���XiE�Lr*����a��<��4ҧ��%e�zL˧����CC�E�?c��R �pj��;|��Nz O����l�Y�0��Q��2Z:������~���B>��ĳș3O?�f*��R���Y`�7�������#�`8ā�-,ho� ������^)��u��pkf^U���Sk"|els$�ޛ����+�ͼ�����CP}�]�K�,��qH��v�>�h�q�N�|�Y�%u�e4�����~ZL��Z���Gɺ��.ET?��_�����0����g��ر���������m�WqT�V]��u\43�	� �K	u���G� b&�F��+�: �| �	�u��I~HT"���{�J�6T�k@6����y���D�S�Y#2�)�Vpk����'f��K������rҜqLo��h���$EY���u�f�t�O�?I����'ȝ'���6��l��#Y��RZ�{�a�T9Tg>e��у�T��M�>��$-;�[;�ix^k��f�`���F���w6�X����A���#�}J�m�9���lZT�nS�#+����.URt����>�����u���c)M�]�Mr�H|Wa�Þ_&-���JlЉ&�KnQ ��C�B�t �}��Ƀ �#�����u��1m�||<͡���r+��Y��V��3O�[��)=�<���I���Z�S�ޭ	8U��O"�t���c����M���#<�>l�+R����@�z�j.��y��2��=�Uͨ����O�U*j�9��a|f|pN��܎��?��1b�IM���T��Y:(|\�u8L�4΁6VT��y��8X<��5;B�mN�5��\+����tsҚ�e���ʑEp�Wۺ��Cu����x&M���D���S��y�+� �7��,�*6���<�W���qB��·P��^�s(�?9-xC�)���K�d��{Y<u�����"m����.)	�ەe	��� G� :
Ê��	�"�E�uF�4�D_{S :�Xo����C���E%�L2�ƒ�;F�
��!���U�����)t�>���i�:�t���[�9-g�pU�d�|��QwIH��8��Su�}m��m����&RȽ�f���X5�<F���>��[�ý�������%D������ QA�և��)]yz��[���"��Bea,�9G�J�qT�I�`��ѓ�!����]�>
��z{��S5�#;s�Ў���.n�&U�CQ(���cOK�u ���n2I���ǋ}OE�V�S���ר:kgC�0�ݡl�b
��Q��w�0��@R�p�C�/�A�<��#�[]�M��J�υ��.4�q�F<"�1�
tL��
d���_1^�
�iG{�ֳ�[LHO�rW�G3g^�����pd`V!~���1��cb`�-
 ;�2�mf��dqS�3O�ӵ�h�|�.hh'��<���P�h0���v�
u��2OK��9|]X�0Ƞ��W�l��Ֆ&h���_DT����6�8�������*��·5�y����	K]�;R�;dL��W��&jCΌK�/׈��:�bA�N=�:�AZ]���1w��B��ɜ�}P�B+�D� ܣz;�	����qD3K��{/}�0��$	�@��y�d�EU3���v9���4a��b�G�vs�d��}s��:j�>w�=[!1�ulc��;���<	֝>�0�t!�����P�[��O<�ء@����� M���Ti�"Be�e6NE#�.}>3��Z���* T*�"C�&�6�Y�<����^[�oӵ���ט�:��Vj9�Q0��&�a�uD�>-���9e�4U;����U��ᕴ�|����ʫ�X���>9�_ʅ|�!sb�T�AEiB]r��5���7���)R9c$�x�o�#yi�F,v���-jb�BZBZ^}��i�i1��R��A��n�9'5<��_)3�m�%�J���3��{dS�k�eF�yw�V��L�sr�i��Z�%o���qV<*]q��v9� ��<ǰ�+)P()�hgmG��%�.;D�Bh(BS��
��/�7E{ܐ&���q�_L�O�;�I��F$lн	H�
�S��	}`�t� ��S��u�l{�F�sS��R������4oz���[7��	���TO?��/��r��W9w;6ܚn>b�m��=t�j�1��FF�� FӀ�_8ẍ́�A���ȴd
FM���6S�/[7�� U�_�)��eG�תyE�<�9�F5����l�X��S`Ѐw�~�l ��4�/
��Q-=R�� G��>ޗU^�����z�C;��PG2�����h��4�s]�e�k��R�(��g�\9��w�ݖ3	��ҁ�2WBo��e}叡��S~���N��egJ�ǋHeT2 8�K�{E~\���]JMR�[t���g�^ }�OL���/��p�s�� ���%|�aM�dX��2��@����P��IHR�2�ʬx%1hđ�ʊ��;9mx}_i�ω6���*�*9S��ȕ���B��t�d�Q�k�-n���A�Me��������n������9��v���"�e\~=�ߦ��^�����o�����{��G:�Uɿא� }�yc�2
kxw�D���ǉ̹c]�9���9���mbũ��U�]S3%'����cc/Ӊޏ#� @����c�8J�X�F���֟����*?0�Y��!��?f�0�4x��5�f�/A[}�/���_'<�V��c&�y^Ʌ�5,j�+�o�����ƻ�U���$�7pᮚL�Oz�V��+��t���G�T��.��.p�,Z�����V	���d����i��'�qG�_�w����8jU�,h��EG��-'�������F������=�Wݾ�2�W�b�t|�fz���_ŵ�UzR4��R���>g܎֫���V�w����I7[�{�]�Y��s�[5������L���2�e2�%�)����C�*��k���[�ӊe��n�������[�W~��䨉���݁د��T�vN.n�G�90�2> d]�w�p�a��+���:	�bl���	(\���:�^9We��h���'���@�p&�`D���:����� ����Qk_��<�h�ͥZCm�'�x��BPy�m���B��q`������g��^m�pP2)���#K4jo���B1fcCB\��S[�8e�R�+�"El�!��D��P��-���ɎڷM���a�BzA������ R@�sB�u%H����G��L�N/�8���V�-�(���N����8�*z}��ά�&7��:v҉J����"�U�v9�#�*��јT�'�Q��T�l軙���h,3��D!Jel��o_e|���a/\�5 ��#��^y��葬��>I/�J�-E�^e	���[��DĚ��#Ɋ��Dh��ach�ʵN��pYc��-Kh�*���x�"�-�l���&]��/�˜�7���ɿ��+�Q8�U�q36?nWNjr"M�e�?/���ϧ����a;x.�㩎<$����/ǧ(晞�0���������GFi�\�݌m�oz�YlX��『��y՘�=w5�4�:�� ]�.]�<�΄�-�s.�ЬE�pV�k�U�t��G���n&O���@gr�N��C`���{��}a�4s��6=ʪխ�ݽ�I0�\mГ7�B�G&������m��5_��1<:؇�i���$��e��Z�@�$��/��a��t����a%CrB&��{�8���-�����D����C��rc��YY�5D�=9��Tce�k݀�#� �%�1���ͫ�tg��G:č��d�!����������/hMh%��Mɐ�:�.���
�'�yԏ8 '
����Y[�P�8rD�l��~�7���1�y�f��%�"$?� uR��#w��M��Ѣ�@{��7���I/��������n`"�9��GЅ?����xZ��^����ML�wh�m�xX�ݞ��H���� ��k���<���OVm�/�S�)���Fa�>���. �=�aX�=�Y�W�tR?'����V���HN��μ�x�_�ͽ���uR��1�Dl��",=`"�����	�V�OX-a���h��6�M5!�dU��V��	.�5�rm���5���?� |]s#��� �-�c��B���Yg{��(/�bO��|��-����|�D�K��<P��*rd{���(i��`*`T;D���p���}�	~ ������A����U��΢�wq�a�G���Џ����#�d3,n� @F�-��`m������(�u��,�r�_���ox��A�L�VD#�Z'���ܤb>���<,�����f!��Qb4N�b�!|�:�.��[ k5wN!�TE�/���E
1+p��M�����J��]M:>��VP�M �tx?��x=NKR����%־�3PNƁj���"2���2?k���wS-�[yM���z���DEHZGv��DK��
CKM�t]LRy��n@}��
�Go�djњZ�x��gM�\o��G}�����I��{���K
�=&�i�����r�@����c�ш�����i�'hi
y�0���k���T�#�cw��>! X.��q'��_��:�ē��$��eDz��Th�-G�s��ϸ��P�[9�V��� ��l��8����}I�C�P��X[u}���o��٠[gp赇r���HE��uN9z�؁�-x~QZ������402���1c��c�],L'�Y�W�RK��-"cj�J󹏵��?:H�0��v��ϵ�F��2Uyn�&Te��EtB��Y·?0���HH<5�&%�L�]�)���v��aaJ�_�W��.F)��%d��d��Jh$C�:'�'�?W�5�Pca�;�/Ȕ��lH)� "P󐲤�hB�&!�B�]��O�S�0T�_�~jǢ"�~lR>�ϐ��6|S�c~�@��u�li6g<t�R<No����r�b��4۰Lx,�!���^�N,��Dߞ��Q�W�9r�L!6� ��$�ڒO������%3�$� ɾ����C�ڭ.ë�y�ΐ����5Ą����#9�ZQ���V���f����I6���ڈ���)��(�{vb�U��%Z�����^�]B���OQ������xB+��<�H�6A!SG���u�KD�+�뼀����$N��)�@��{>�K�Es:���:!3�|�F����D���>ҭӟ�i���|��X��4��~��#�ۿ��A`S,�	x���i،G��� L&U�B�u2�J4Lwa@?�8���a�ԇ�B�h�#a�,��j�'k�l�L��n���S+}T��X7�`���;7,��ъ���ErjC2.�3իP!���iO8��ot��S�A��žOPa#m�
J�!1/���=��$@���@�2d�Bs��Q�Ie �	������ ���t�f!�i �n��MR���S��<K �j�x���:�=����`:(x�
cCQ�U�L�[aaDK�qN�����Q��rkf^׵��-ϘS�)	`'7Qpg�ʝy�8=�8� |=
� ���|#�ߦv�\��D��8�ec�/w魣��O3����i}��&^�>�~��3��U�]0����pY&Fq����S_�t��0)��EV�?��S�����{g���%�[�cp�lɩ��Q�����V�:�򱈲%��.��t9�Z�icڸU�VeAe'^SP4�����,¤qf�"���k^����C��5	�y�AB���P!��	gfU�+Ј�����3�nPPc�Eq��)P<b���e5$y�/��x��1_�H�'`��߿8�o��i���/58#n�sR����3��X��XMU�/�@}{V;�۩�;�r�KNZz�y3�)�I������p���-�)���ӑ̤Ȯ�֍�@k����[F�'��UJ� �A;I� ��@��eR�����S#[L�tx�P����d[gn��b.dk�R颜�Z��
QKp�T^|x
i+w��d5����`E$�^N-g��:)��R�{m,h�k�`Xʥ;��K��m�t1�����U�d�1�g8J�*�*:�k1� �~5��]����m��I��c�P�ӖzN��m�k�	��|���ڣFf����jX;�W�{��r$�ߍ*�Ew�y��
�<����[��xu�+���Y�(�7�W��Cc��ϔ�Cz8���~z�!z��g~�n�<k��罁eZ.6��0�X̟�?��_�@�{�t�	 ا�!H_�Џ6DUU0ګZf?�)�=!s�L�	��1���_$�&/�'�@{
��g��S���H�j��Y�H��� Fq|�70��Y��w�ȧ���K.�lm��=A
�fĸ	��T�f��FF��n8��X˩�>8�!�B]_�����2�_ yzy@��@�(��H�X�*]�}좃ߌ�.�&�/Ѐ��Ŷ�����4�����i�=g�F԰��#��r�h_�9˱:R}�=�	(o2&�����(BRSF���p�ϔǗ\�Ÿ�J� ���`yxOLi�X���j}�Q8H;X��>���]b1-E:�m>b_1	��W �fu��R�$���d�eC�ٟ[�j ����gOzLp����:�Ck!�3>�F��$�is=��;���I1A�p����Wc�?�j�����W�{��=p�L������v�T���S��.��ڵn�Æ�$wd�+!)��.��EǏ~��e���4Ff����^�,x7�)4��X���7>�$�Y�>W�J��Q]C`kc;	-�H����ϭ��d���}I�Ѕ���T� ?ld�%�V�)��/�l��Tᴏ���	�XOad͜vh���-�j�d��|�4$C���#����G�"��e�-��Je:���������R("����Fѯ� �$/�<�ۛ'�����ùf)@э�]����䃁s��@����X���=�+���ZD�@@�Dy�ٟ9�)6񚽅����^XK�yq�'���Z�� �`�[T�8B�/��������ح��&�`��ZE���X"�������3[�r9ێW["�n��߸�퇄��u�-��CTH鑺oD���~W@�V�\�Z1�#�F���mm������\f� �̑q���^�y!\�<R��d����Z&�q#%���k��t�Pm_s�>�{җ	����zR��a;��k�o���-sS���L^�vx�����Jj*~_?�l`j�7��_�����/n�K��}L4$,EZ��o`4.q�pƏ��m����Pik����{W
zC�K�����u�W������̿z^�;�Z���*�����}IЏ0�fȉw��}0�����Vwt�d�J������_�[���o��a�p�x��K�|�z������*��vP��\8�,/�����_U^�+*���P�.�����VEd�l ����w���y����Y�T�ؠ�E�!L�ȐV���,4�U�Y9��Wr^�)�oAA?�Ѩqz�,��4r��s=	5�;�K�K�_[�	���U�F�w(�5iO�4ckF�r��Su�*=�����Xέ���_��� �9u�������_2�#2��E��~X0�)Z�?�V	,�m����,��ЄJ����
�[f�v^����|d|Gf�q�|J3�s��cy�[��RW�}/H2It.K��6f��ؿ�v�}}�~���0��\�y�?w��s�
W�@-��Mj_�&4\4ɬ^E1՘�y�qR�3�}L�P��wm=.�Mċ��E��z��N{�a�a�Zh�����ֿ�"�G�/��(W�O�ŵb�\hU��G�Q��:i^0y!2Q>l�0P���T���쒒J{���\+�����d?͇w-��`�Lٜ4����*o������h5&e���=a��<��(�BBH�#�����d���_2��1�=��ƪ���k��~! �'$���\��=�|�N���J�{��%�
9�.~� ;�J���*�\MV1�]^�ÿ́�I�HW�$brOc]�^}U���v�6n�h�%YF�LѿE����0���Y��-m[�!%�f�z�@����*4j��Ur;{Hmؕ�Qc��(k�T,6���cy��Ei$���������y�Et
��-cK�߆m(����<��kߗE�����S��ːf��P{so}Cz�Ȇ�夓|�� %�ols�A��#p���{��! ��|�́:���ɲ5���y�@6ʑl1���u�]�P Ve|��oE�to0ư�w�8ށ�v��A�;Ot{P�v]���Qr��oLY�hI6,^��A�妥�ծ��~n��A=i��y���Ce���l�l��:�]��`<.�[���t ���Tc��L
	�s�Ru����՟=:{IFc��e���x���|Ge�w��>=�SA��+W	�.8�� D����[u�%��H۴��7ɺͦҝ��-��_��/�����CV��I�q���݌s�����|0��f��[d+V��Zn��r�^gj]����ڏԖ>v���d��)�_H>Ң[��5�S���g�B\5���\U&�Yh�)��V�A�˸_52�DN��|���@�.��6*��wzrd��H;���k��˸}�����q!@�;����
IDAE���r��BZL�8�/����e�l�X�4_�V�3a�ސ>�.��&qz�^�+t�,h��J�6������R��Hn6i��������>- ���dˉ��m��q�ܚy��a���3ܕ.ޙr�jl�L7"qSĦ�mե{�o��N�<��n�.�<
�	w0�gs��.�O�,u��z��fڵDUV'?܂.���EA$���7�]���R��g��;˚���2u�].���%n^�X�����J7ב!1Q�U<;�ZX�i���8�{E"�n�ꂞ;(��\�7���H:�wA�|�g`���՝.��xȉi5�y�"�VQ �r�W���<��xt�{��M�QJfۘ�d�HZ���#��$�̟*6�auZٟ%Dӱ)=;�`V��=�5x"�d�����q�Ν	oW����(���M���y�:���X�6��?LOPA!�����B�R�o�a81%���f,E�phRlO�Yx�e�X���=���}�M~e��^��G�&i��N� �y�w6hE��2����2� f;u�iiey�"�N���E	�*I�z���j��p6|�K�>P:T��a��믴Zz��S� ��=C�Y�5�R��l��w���B��6� �]2ͫ������9b�y͗#�p(~�Y\��:���@)`gr��.���f&��!L,�<��`��~�ʇ���:�f@��YY7ܶ�E��\�Wu��O��2Th�*jk��,�O��e�t�K��-�H��n5���C?���K�t��L]�|n�4��P��_\��mͶ���yड़4��~I�+�#��M:3�a�gS3\J~F�C��hHgC/`�Ү� )�/�*�`���ggR��ك��RDf���1;o����K�=��Cz��g��0I7�pU�r�!f�R���	3�>�W=<�K�	l;�P<D���͆�M��CC��
�p��9��7�X��y 1���)d
l�&⟖��:#Ɖ=��>G�&�3������X�M���nUV�*]���c>��B�#\'-��z��̵z�B����lq� W�=�a��~�oC�AQ��\��-��Ґ���#�eӀ��ɩ�(ÞW���3��^3T��u1�n��=��d\^`Р��`7��:�nL��:J��Ğӫh��?'q��Ԫk���Vv���4���/����-�i:5~iD��2E6��7{��䌝�du��)^�,��o:��
@����Lq�l�,��a^vu/Jnt��_�1ߔ�,d�{ב{N����{:�ȡM��ߦo�E̪w?�-�㱅\�M\��蝥�鷖�v+eɢ����c����U]�M�n^f�:G��6䭮�9؍�(p��T�\�w|zt��(0IEZ�����L�[�l���RA[�Tt�q��	���l�k�'���_e�?Y2=��><�M�R�;&[Jl΄[��I�?��(�%s��z�I��5��׈X]rr1�m�G+Po7�=���s5::n�/�����g9Q�F��Ed�p�Ŕ;4��4ǹ��PZ�[�
�2���Ů��~PՈ��<��T`�,�$<�@�9���~�?5�g|�`ZºzH���	f��S8ԁ:���͘��S��u��a`oP��p1]�Ϧ1��U��8�R��}����>�Plq�h�;'m�����Urr�~��Z����W��;k�"��g��@M��"��
���>%\�`�o?ߖ�-��f�W�|Kh�Q��(��$Ɲ�	��C
g�|q��)�!��I>��~Kñ���;(*���=Bځ�|˭���h������_T<��*�ހ�#�y�u;����'����|*5��}֓���v���X9��J�.�c#v�W�+��Ua�{�&���O��ټ`L+Y�w�T_�,�_��7I�������D