��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U����*��1�n<��V����I�0=<�i\�	®���PDo��?�3f���E��!�eYK�b=���ؗ�������%�0�#��?�	�Ol�ST��0
�p>�9�^�ɶ�V����ba$����~0�^aӰwN��S���O´�}����`����C�h�i>><�H�ھ����`�լo��Gn]O���=a�o��V8$�l��:|K0"1xqư�';gmC�����b�]4>`��|2�3�Z�:b����M��/�.�A}��aW��q�2&�QtkU)7�~��%A-ߎ�w��\i�L����A��X������D
���.ފuoo����mӈvv����N�#jQ���H"��F���eׂe��n�P0vw���.��W�)+�6�8�j0�D��D[�ʉ�V޵؃e�;k�������s[o�>��a�Q��z�y�JG5�	Oֈ�=M��E�h�r)�Hz��-�
?g���7����v�>lFa.Q-���mN�]L��`~HDx�C踝;Ep;�`<c���>�ُJ�iݮ�����&�߷��]��BF>^��h��̾�P
�	E��
�m�h�|��W6
���Õ)�����
��&Ƈ8p�_�y_�k���K���>�Ph9;^��aI_�N���R����-�Ӂq	�:�S�va���&l��"}R����v"���!�c��=��%>�}�c�mQa�ZE&{�6z��Ts�����C��p���u��p��-�٫�-#Bn
t<��6`޵ʈ5�O��T=�����k������P	�O> M�V@^��ea7�����S��^9��_s/8PL�5�w�� ��#j[G�o��;�Dz�K"�]�#;u;��s&Ӭ�/�s*U�U�%����e�m��l��
Ƕ������[�G��!d�db<�F0ٚٯc�'�,��?�LL��
�F��;(�&�~Tm��R/�v�T�"���PÖ\�-�O�X�y������~�tC��S���t�X��@n�4qn�� ����ȝ�Cp��	Z&�����L�d�tqﲄZ1I��8���$*��B2�ܢE���t��VtT�]�8�9����]�\�a�p�D�Qh���bV��T��[�*��ULX$H3��l�T�][K#������$���ʿZZ���8(g2�s>�	�(e�:���ƺ:����gN1�xgE��ebK���[zலف�A ���	�|��e�y�W3~x1�/�L��������O.��`	�#���*�0��q��& *�3+����;��3.&sI��1~���\�`q�%F+Y��a�b@tc{o�@����"s�@~�S�r*"afL�`6�U�����aQ��X�B `�M}4�Č>� v�K�հAիݚ���}�5����|͋�j`ª�0�%��I�3
��/J����P��Kŗ��]���-].�"#)�'h�k;L��_�A�q�U')��QIGd�3��z���.F;�����_�D�(�M
�H[$��B��G]7(�e�d$؞x6�`h@o6\v��pvpE�o��*P�� l)���/Kƴ����l���<pPv�1��)�b3��U�F�Ι5a����qE���02�s����l��X��6���2�-��{N6h޶���æR<��Mi�(��}׶�V�8�&..0�JQM6�����Ԏ�BF��@R�>��d���2���������aǟ�a�V�V]�F\I.r�M��N��q_  ,��[�U����PX�_�_��T�XVOcX�
K�3��Ҳ�f�{��tC6��ȱ�f.:�^=�#R�`���r�嘳���@�����uhҋ�ؿ6X�� ��1q#վF����F�3h�o��0;������~�����/@o�l\Z�$�:J�-�����R8H!�)2�� !=BPx���~�g6@Y���gK{���	��s���� 5�O�Uk$*�FS���]�����WI��%��9_��"[=Z���+V�EV���iVY�R��m�8D;KB.p�~��Ol�Q|yr0����,9�2?�m��i�US�P#�'Q�	PQ"`�0�?��V�MZ�dX�z�˃;R���������V]��������с� �]b��C<�E�\�1��2�J�<�8S������0��?�� >�c���/ڥ�Z���i>U=�Ą	�8*��]El�4/�)���9��Q�=�J�>ݬxv�鸹����{�� ��eʊ$��8��q!x��7��S�)=����k��ܡ��g�����sL��K1���+���{җ�e��|�b����x�.?���W�#%5�Բ��[0
��M6�tۺ���AN+ ��u�U� �{)ߓ'L&���u�	�"t-y��w3��b^�����Y��
H���4�l_K�ʈHA�S{��d��ŷ��$����}�I��4��|����1�A+��^�LW�`�k��\�x4��}#�Í��g�Φ*���
h��@���~��Yoy#&����/̬Ĳ޼&c��9��oa)�|�OB�1;"6��V���Ey������������|��u~_1G���Z��J_�n�Zkp�]�� {c���!�L{C/o���'��T��Լro�2X�s�4���v�8�?�����kR*g����Ą��.2]�ݽ}VdB�����&䟹NE���������<�G�Z�7�hq|_���f���������\݄\�$�*�+4��1�ǁ@���yt���?_��SR�°U�� ��i�)�;gz��?�Mk6A���hwT^&I����_���CX�F+�\Q_0���>��C��}y�l|�������5�M�

o��ZQ`�3=\���<���*9YH��ɢ�����qѿb��Yʝ���mP{ʻ� �:^�m!�w`݀�tF�����z0�3�j�3�S�bݎ�?���F�ls�{�mw���nձ��C`��pe��z�,M/}fZDܟn�T�?%U������(*3����s���LT���a�4��HhQ|
g�F1����ӱ�^�s:.J�{M  ��϶�3��['θ��W�8\ �|�`{e�"ѿ���:��9k9�^Q�E����Up��.�w+��a�z(L�%8�D)Y-/k^Z�r@S8J�D�V�C<���h�e�'$���(DM(>A�x�w��m��`�J1���p�Mw�b7�oÀ(�S�x���P�̗�X:��ܐ�7��º�~�Th9�nZI�͉ �f�4�6�x�F�V�.S#�q�}�S�9�(��z�;Б������#���M���^��!ݩ/�J���/�/����42g����"�L)R�Ɵ�éwr+$��-iO!��m�r`�q����-JM��?�8�hJ��� �{�"X�GH�����U�PJ9@���)��2�����k��hH����Ԋ�S�S�)�c�%p�p)�x�hf��}�D&�؞2r��BV���U��Lf���k/�g'��jRX#w����d�������
���6����j��>�h�Qx�V^�3/F��$��V�R_��o��\�O�%�'�}�z���f��q$p[rE��!G�����.�F��B�6�G-1q_��v\)"��;�}h����̤��T7@�3��]�H"&���$1�p�?���0���5yJw}<{A*S�[�{1::e�� ���������a��z3x�4��8�XI��ʖ3����V��l�q�bR���x�_]�,���ԋ��
�/>\0�kV�v��~1V�����@+�(�}�X��O���y�T�$(��ڔ��@��RN�K���7��w��A�*��8���*P^��ˏ"��z���}*.~��~h��4�R5��T���Nӕ~S�x��:D*[:5�Q[�yŽY20�
�#�+�W�5�^ 	��W��J�(!���(i��ȕ;X���Aؙ]�Y��z�&�
2-�\�";��S��a���<�}띍J�ۄ{���R�,�v۩�
�4N�3�&�q[]B٢ahm����n�O芳z���H��Hu�P������Tl�#*����$gօ࿀�[���Ί8�GH!���f�˺�Zv i�����ԥ���#����\E�j��xK�2��8"HuD��gc�^p!�l��ᗶ�CGDF�mu�-�����=�`�<��sX` ~{o��f�)�E�6|�3��E�f�Ln8�$mϣr���ۉ�n��B[iF����~>˓B�dQ"u�N����"�N�A��^�v��բ�|k�3�L�dU�j��?)� 0�d�YGwF��靥�z'y�}ey�䀏	�Z�Q�}���C�&Z��N�@�ǫ^5����n�-���M
�]�R��d
ou%Km+y�����"�gn^!x�����`�˪Q���}*�3��k/ox!�7�M����}��vѣn͆[���QP�~���꜉����Q+|�%��[��~~/��������F�~)V?�R�˟�`�:;b��;*#/�\����Vo(��"���<5��h�GRJq���`r���_/y�56����M>Yg����Ća��)�vG���
���l?���ocC��]"���v��g��M�0c�g���e�۸0k�{���46޳D����˹qA���Xm��A^� "&�}9a2��j
s�;9��$��h)o�"nlx�8qǍE}W/̪y�nN�כ���R���$�>` ��n' P��k��'���L譤~Y:�����+�y�Q?L��K��&C'l{�����V�����s/�|iPb�`�8�*9��C�R]��l�F�&[�.:N�!�Z[���u��T!��QD+#v�d%L�{Th�CWy:�������ԯN��ݒ����9��L�8H2V!w��^'��K�p�3�@� ����WL�iz��殕��F~F��J�$�HK��F��"R1^�ٶ*Mf�*v�~�N���ex� ��'��{0�e���m��y��5U+˔x��
��yp|9 ��3��RK���.���_��{�N��B̛ɫ(*?��옊u$jk\k �/[�Jb{� �i��,i�������m�/���D���XKR���Y�*(�np���J����E�%��@�=�������z)A�҅�&^�ʧ@p���.`�s�~��:�ٰ��nx��bଊq��s���e�\���a���jv�hd'�	��$��9r_�x�uUG���0��N�f��?Ƃن��?���-S/�J�VM����F]�	|g^^İ��V/��Q�k��*��xu�
�>�[�l>�9P�b�"�=�D��9�IQ��%��E�%B�qˇf[D
ȭCBj�8?��I�	���\
��|��|d}\&w�i�Dfc���U)׺�DM�vJ�ē��?��2>H#�E�eTr�)��D#���ܢ�hok������'��ݜ����|Eb~�3/􁧳����g��4���t� |!�eY��5��2���?��� �����W�h����N�������̄���c�������d����_��&�c�S�:^��S�C��;T9O�H�IE�����~V,^�RU�R�n鈺��n� c��Y�y��8���jm�$�5����ݐ3	�nY�����`��O5�()(��-;��Z�������huowz��������Z+���s�	�B��n?��!ȤzZǊ�e����X�C�����tjK����@+�1z}ދ(�2�d�W\i�lg�
ܡ�]�{���%p�yU���"nO���f�s��vv-[\��Bjʙ��ܡ�tOcknt:L���K&8A#��j�>c��̫��
��	��v�ܙ��TMu5�y
�욹Ϥ\���!�?)�9c@�/M)Jl� kyhtĐ�DI��򍘬�a~�I >խ�hP��*�WL���rй�
��h�H����W���1{RCVCő�"���I�,Y�s˯���]��e���z�Sn��De�:H��<��}f�6�=�_n�8n��W��ـ��B�YD(Z4q�mli�pg5b~�H~!:�Rb?QAG���I�FP��^�'a���w�ܼ�n�@bS-Li��e�Q\	�d��-�`衑�ʨ���0�<�^�xo��~5�nJ�,	_�o�=�os��uJͦ�(�O�3;t�g���+rl��_>�N��Ϝ���D�s��_%�V!��o��zULd Jb;�f�Z��� �/i��Z��M��M�}�ˀ��ʗ�3F�]5(m��}n�u�� {�&�ɂL��ݒ��M�@hY�;��.b�����[�n
���t�T0*K��օ.�we���>H�"p0. ��uw��l@E{��bm�}�N��%���r���V���9C>�x�h�!�� ��$0��Բ�6��� ��SHL��b{��Pb7����X��N���`�B�Z;�7�� 8��� �b	�/~��*)MXe��T�L�$�{���מ�ń �]*��W�����������kaP�<���Ff9����+�9��Yc&r@���O~���Jݖ��*_?z����z4��m��*DZ�5�ЋY�H�zt��%�C�,�?b�Hhy�g5�X�C |����YMK�-쉭i��88�`�!5
�mV	���Hg�pd�#�}��p+'�C�KJQ��S��(���[{���GYU�K����sg���gq�����ijkn@����c��~��ㄧ��M�#G;�|�1��z����KB䔟�?P�F
�bk����
��za�(�H���V�:
6``A��=�"\`���BX�P��(�.��2�I���/�]-��O�ݱQ��҅`2��{�CU�pTJ넲d�d���q��$�[����L �+�'�� ^�VF$�FY⩲ۚV����U8ʂ�WԠ����sԦ�	G��ib��*��an
�u����w��zbA��L�tFtۆ���fo|2�_���6(��S�1���d�C�l���&�~�_���B���ۜ�љG��z�`�9W'X��~y��b
���"��;g�*�j���f�e�Q�F*I9���!u� 5��p/� ���yi;�GAe9�{0o.<��ɩʸ���:�)��[�0��l��)<��.��]������ź�|S.DM&��rvǼA�c����� u��t~�?�2�MV½�E����д�e(�m��Tq1�A��i��A��|o�_���u� #�s���JOX`�N�7{ܒ#����A�d~Q<���dSŒ�	�O0�����ʦ�~c�qL��/�f��M���z��f�� ��_=^e�oQ�m�OǼK��)Xt��/�υn��'��4,�M��ޑYq�+O���P�f��P����ǝ���F��2�4)sū% �6�1��Q�G��V���U=8���x�^G*RK��B�3��:6.O6���XB�ĭϝҺ�I���NE�S�Y�t��!�P?*;E�b����f���-N'7�X]F�h�u�Wt���J���y�N�5����i�e��DY��Pv=O�b�Q|�굿�P����%���j@W��Lj����(J@�b�k��3S3��I�,Y�� ��ѐ�-�nT#n#o�Ð�f��fmt�mв���ߐ�M�qx!���9�d\���r�������W3K��qD�@��W�<�g'O0�2�Vz����W]�&i�/vCڐ��W�ɹZ�LX��w��;j"_Cux��[Y�:��� �\J�Ÿ*'{>v��N���߱.��s����G���h
��E� ={OB�l�4��#����<���'d��4�w yt�ق�d�J���{@��]Ty5�z�D�o�&��W�(����0��n3����@v����ў���Z�:h��R7ߝ��D��X6,h<�Z���?�֒�c|`��+lO��
 s Gl)o�2�$�*��*��ݚ�a\�ɰ�M��N&Kw��h��@`��DE��Q���4cH��j(�a�LC\�SY'��Z�J���fc�1�9#�Y�̏4,��j\�����N�T�Ny��lQ aė�R�5�܌��;?3�'_gD[�*R���,�|�L���ޯԺ�4;,f���\���+ߜQ5̬\�a��;��_>}�����9uK�?�w���A���Z�uk�&���GEbj�SEd������^��<�xN�� f^�P�{��&�o�`�tm_yLV*��p��Cel�!#�^���5b�c��Y
��K�&��B��`Y|�4���Ư�!'���L���|���pe������A}�y��ul�