��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��¿�8/�L7����#^<x~��=Mϑ?��F�D�H�:���3J` �>����e�|����*����%Dqa���G"o��]6n?��n3�v�{[Dg|ƁP0�JF���(��@�w�-A��zF�����<l������Ca�r������T��q�d�l9szuB���O�	"�Qj&�y��9�PH�h�R�.�G�Բ�*��l��p���6��A��|���^�'70��0u��$�>�F߲�,�Õ�pS�~j���]_��T�N�\�p�1t����Q��.�����Z����[���NF�G>��/}�����P�%e��'*I���Y�x�%�Aj����	��J:���|��
�������C���6���9��bRZJ�@�ڡ�K_j� ѩ��%���z��d�PA�[����14r��U���@��/ɵFc�zX���̖PKg�Sl��ޝ6�j���Yn2��C����Tq���a�T�J��ߏ��BF�.�dD��uO������X��Yɦ0�'hF
�q8o�D�-{��8�`��}�<r�w�Z�uY4�V�@�v���o�����TG��� �%��ҳg�O�v�����Y�ky�/k%����~~�};�a��W78~W͈�i��z!umC��5#Ј����ͱ�,�)�0����=�?��;^���7����J�.E��\��N����{� �Y�Վ�#��\4�Sc�X���w[�HpJ;w��O�(�6��3�9��^+��|�j�L��@N�Z���m�1ђ�KI�:�+.�[��C���k����b3��Zu�y���>S��6^q(L��,$b��>u����#�)�Tݿ�,���~F~�:���Z=��5z:��_��6P=Һ~��@L_)]�����`�����@��eI��h��(�+�.��t2�#ݣ^��N���3U����\�$T�=��}�zV��&�awm �o�����t��4grNR��Cqn�vv8��8���@��"2�hY�R*Z�&�v^QEtD��!.��cѭ�_�n,"�us>(�3t��MF��N��1'����/��
*����5#ԡ�;8.��Xэ���	Jjg���Xzϡ���$�� �w�nˏO9����Ԃ�î�|M0�o�F5��o!�*(#�u淎� �<�������|��U^�= �__t`���O��Udu��Ȯ��1w'�$�9�=� �{��^�*$-�n��ɬU��W����3��/�o�3V��2��h�_ƳdD��Sp���O؍�]V�!�;\٣�����m�4�~1��L����x3�wO;+�MET�Zu�#����@?�/p#�����)SL@�Dy��a��h:�=��
)� B/՘���Wl�P+�z���63�N_`F&���҆h_(�\��� �����2�V��<p�G� G�7��:��`�X���$�&ΪY�Lk~*�zL#�gM!:�Bj�����+]��:I�Cd5��S�#MH8uL�	")��=}v�6:
��37�>��@} ��	b Cu:�>�v7�^J�o��K\/Cx���_9�p�Ҋd��^�.6�f�:.wBz��#/�怵-���?�7�ƻI����:�"�%�V�S0��\z̫�\$�
���c�ls�D�tZ���n�l��x��z����wfp!�������x
�y���������@h��C\�I�ΔV�٥�ZS;�Q=��>/���<��`��!-�ا�y��{���2���>�A�t�X�?��_ �
��<�QK���$�b�aß�|١T���W`Ǡ�.�~abf
��"�oY�B6w�t7�\�:Gc�{����S�@�{F��T��{�D
�����._��?p��GcD]����퍗�U�*��L��Ҝ��f��՘\�)]̇V`�c�p���f��2\�=>A��:W�P���C��x�G)�~����H�f`��Km�l�f���&��J��wU�O�D%�W���9*f�4� '&�d�XX�>��8'��hTJ����|��$����@����i��Z���Q����Z�hyy&�Ǡ����CzB���vH�9�)^S�jd	��7
��L"���t����G��ݜ|i�� ʀ%z*��Y�
g���>������Yѳ�N�?z$�
�?X�ͫBW��|tf�'�{><Kc
����B�|gW��oJ�a��\����jg�*�=ٰ{���$�4JMu�<`���q���3m}�8hOo��t"6��ƦMh��n�')E΢��$�=�V0F#*WC|.�]��>L�uS�?��J��T6��?5.^��1MQe\���Z�"{��
6�P�A
c_(��9@N�>�i�
nٵ�a�=!�B���*��i}e�g��E�r���:�	%�a�;��j�'��i��k��0;�ܜs����E�����Q槏����(Շe�x)�S�#�u@���$nʙ�T�Gu�0���`��W�債��^i#RC��X���k��Wc��&�
���nV�;�x=���m(��C�ylv=�
�O;M����[&��W#���T�m$���e�����}/������8�*�L�0ogߚ�#�;�s�ѓ��|t��{�o"U�G����;�J�"�HS��7��,7���9�4���Pw�{� ��kF)~J����!�o���������}�W�>�&e���?1J�-�0�����8اn>�v�D��N�C���������D��z��FiWs�j�����\Z��ɤW��㶸�8_T��5�h �Ž�<(��K�-N�7�K�(�FG`��%�3�=:�����@�KHAl��H ��f�f������vy���C�83B�zz�B4��AL#k�HذH��P٤�J|!�6+���d^W���{�	�Er�Vȓ��\6p�`��1;��3PC�-�6�x�����tQ�3gh���J���dӳ,�i��y]+r�X�7�b�Ͼa����c����`x���
��i:�5�
��=C��+���2��_8�ẟP��k�w*����� ��"Vmg��;�MYh�f?<D�~�8 J��Go*�g��3��\E|"k{�A�ٳ��В��S	��"��[�D!A:$�\ܲ'�Н��g6��FH���3�u� �h�z��^��Vw��ǅ���K�ez�%<FJF�s@ C��d�'J����W\�d@���P�a�xρ2��[�C9F��`���1���>;I�5�&�q���>ѳ,���*e/n��G��!�����#��������/���9g%��Q]׎b�i�+�v�/y����=6��jp�<$�d&���0�"�xzSh����&�Zaن��93�s��	�hbw��ǥ��l)���5O�鿮�7<-J�3�l�'�U�����8�#D��ʜXRT<�D��]ْ�j�M K��r(�j�@n���X%��P?*�$(��pq�]�In,�9k�z�3pz���E&A����E����I	c�x�`X�eQ������n�>;H���t���0�ӑ�Q��cl�Ok��R��D�~GPA	\�P p9���� ]�����jrd:[��q�UQ��o���[Z���OZ��;��V���}�nYC?�f�Ոb5>g�R��ʆ�}�e��t�_� 9�$�/�W����uӜ�+K�K��7�nb /YQ�%W%\�����=����'��ܒ]}��/�_���� �Uޅ�c�
����T�_���rZ=0/"&�
�Al���r*���1�8Z<������p@z����ᗯ�Z�|ʟKK�YÐ�	�ڣ~tk����ڈ����8�}�T$�ז�/� w��	��T�=����^��>�T	���0 ����c^��U��H�!Wvjf���#NPZ?��~��lz�y���ĞS����߽�|Lr/U�7�ҿ B���ɑ&Ţ�m��5)����yD��1�O���+e�T���=��d�,w���n��x��Ru&�6�J���@�'��*���\=\��Q��hk�x��A�=��0+.�� �P���P_�zuG<4��UhZ����lD���C���c�04����g�a%V�a��R�c�|�k.���^cy\�pq���2�C��1��w��E}��s�����k�8Xe�ëϫ���K'�y!���s,0b�t/�و�6��]y���i�4�pɩ@�姃4���Yų:�%0Y� �9��ѭ}l4��w̝�	���N���Kld}�h�We�P��+D/m�z����>���ݜ�1״��*tM:3/�3�:��g�����?/��}8�ة�0��G$���ӭ ������w'I�Q�-)�'��*�EkZ#i����{�\���h��Ru� �2�$5��g1.%�Ř�%��gd��6�Z�ނe�Z�t���+����D�q�X���o`W�?����9�su�������t��j���_�D\G&�YH[���3B�Y����A+e��m��lu��a��kG��;!�P,
��5�:I��b�?Bz�y�;���f�@�hJ�����U�#D�������%�8�1K^)�Hs�ӭ o�9p��:j�{��qP��ߚ �;a�}H�^r��O��I�Ǆw˼��rĹ��׮�k�����7n�<ޚ�{�\#�f� W~�Wt���N��Y6Z {/�m:L�uIP�����9�/��A.J�,������'���� ���*Dgs����a�s��d! �8]��7�&�w�g?�⬋�h&��T�othu�J-�����UGF"�e7%��=
�w�́����P���8�|��ӦN {qmh9��km��P��>�K[�1U��9[������H�t�.᥈7%J�ˢ�f�����v::o�$�H�k��B�T�&�ix�d(���,@b��U&�-�ʰMC��D��"�Ӟ�P�D+��pY/*`7;Ä���������,�Eq��:C�9�T��Ug�I��L��͹Vj�e��>`q��RW�4~C�GWF@���Of���vMF+��u,M��Ϻ���j%�:�':%H������h��;�5����PX%4���k	�.�*���$��8s��&��R17���O�����������Qӛ��1	�"��sOY��"`	f&b������Է��Z%��b �����w��ՒpA����-��c��X�+�C��ϟ"/GI����¬ 5���È5��+q��B�.Ϊ�픣,?pl�7S,j�����`�M�ⅲ�i�X*t�%�[{ȱ�'���Fm�H[Y㬽��j~���Cr����n8E��y�̽�;wr�|b��)�.a?4��l�]��G>��Q&'�v$�x�O�tqTp�Y��w�툊
3 �"�x,|�E4���'>T�Y��F��W��W��U1�Вfdc�0W�&��'��S���c�ؑ���� �=b*DC�[���@zZ8Q�G"{�|�Xﶻq�8�/�{Z��**ϙ��%ޘ'+d	�>}
ޞT��9�!���I\��z�@Q�|&7�v�F����=��NY�\X�E+��$����ͧw2?�DOM �.�Z&�&��ٗ��T��s��;Kf�MI��]j��F&^�n�ϓ���$�9,;4,$��ӟ2�����!�&t���PLt�����B!���G��ho��	�!R!o^z�^�UBq�f�[	ת�	V�q*�Y�ɲ0t�^-A�Iu9�N
|��:���;+����l�{��H3��AV|%ɨ�o�
2�\F �a���uW�1�"R��1P�J=�`i_);�L�}�������I^BƉGu����n�"���NP$����ۤr�p�����F��}����r�9Wu�-6"Ǧ��EL�}b�ټ��[���_�5���?Q����t\�#��L`�#W�^"/mʬ�%P)��'�KX��3�u�*ic:[O�.��V髱����O�	cm	E��*��������}Sy#�;`���s�}6�t+�4�-�*���ض�_\�tT��3h�n��Jp�i��o{ |c���q�-�rH!��D6���W��W����S��#-�p[�g2O�>��>@"�=c�I#�Ԋ�޾ql�=�.�o>)-��e5���3�hwo�t��;Dyj�x�4�g�,;��"/ִ��O�M�w4�VX�n'��=�Gi����ݺ����ȝ�#��S�<y4�ud�BW�V
o��^[���nM�k~�:|g����M^�Óaz���R.���=5�_�2$vX˸��T��^�X�.'	 �R~�S A��P�?�XsR,	���8��lb���s�Oy�xt��Ĩ9�ϲ^ܾ�210ZN�E�K��9�����/�+@(>�4�ZM�2{�����0����vw,�43�ݳ��ohq
��g�di��W��ٔ���0�E�m�q���������R����uJ�泟'ɱ���N��~�S�hx/(��L�X����-(��qs�}���o���� e �sK����)�i8�m���NV�ϙYZޚ+J��v�f4��V�F�I<"^A\Jy�t0�O1��W����;,���;mg���� ��B��:��'�e�`�A�o��TL�J��)w��]2a'�Ԕbw&N���.RD~8�q)������L�1��&����q�5C(������p8y�M�0�GB�༚u�o���4%�!*�;�!RI藖?�
�o�)���-D�ǟ�zI5�{Y��W� YisA�=A�m��@$]�K[��{UV�����4��G[��G"��VY���{�E8�!験�@���Ge�_I�a��k���Y�?Ѡ��xS2�V/����q�kFϖn
~M��V}��z��H��+���Ib9�����\(4�A��V�S���g������NJ�ʜxe�;��Wۋ��8I�=�c�<��0ީ�VZ
4k]���Q�� 
Z~+������bz��a2�v�qR��>���W��o�,(��) ��4�N[/fQk�=�� w�����%D5�!��'���b�Rt����PSZa]n�|�7�fh����N0pNwq�>�[���-%��+��h:��u �o�q2I�Ғ���/ֲ�\i�[��:�폥
��������7���г�A�7�P�ls-�Mz/������a$?, )�{���R���ێ٪N�YD����Ţ��Vd��3�Y>��Ġ��P��e!�Qڦ�w�8b��EZ�i�����)�Cc�&���hKE�Y9$U��R���)q� ��<�ku#f�(�:�/:�������b��`�ܪ�S5ǶԵY��㷱D#+���dڀ��t(�Oc�X�}��z�On������xy�������d.p/2�,����Hx��ҁҳ4�"z�?T[��J��﫚�p�a��T#n�<~�_�|����������(N4Μ�H7�����p�:�~g�h���<M�&8�L�/5R���F��#fu\�5���6S�$�k���ڢ'��|����:�yL��s��7�3��Q񞲀A?r�]'S��M8�"3-�!w{�[^�o>�f�[��F����|+��dJ};�W���d�Z߲&n!�FTĘ����Է,�A�~Dq�ME�	v;w<�1��LE� �`�"|� N����F�eL��J� ���JE��
�m���_�~�x,�@q�Wm��%�kyK٫ب�a����嶥6��:y{NI����b�>�QV���8:���A��0�EI8��K�̌�S��=b�U��lî��Y<Ƴ���g��F�[t�����˽j�z�.ტ��P_�Y���W�5���F1��'�-Aဉ�_�|����f7h^1�Q���g�����ؓ��UJA�*��K���z��`���J0��cG���BY�Ng�U�A��u������J�ܯ���CSn���cP�V+�Z�mp�m>�U��r5#��$t9V+K`�����Fa4��ʢ�P����F��n� ب�"g�l���K��w�8��$Ȥ�s�~5�*�0��lT��$�_�2׵q4)<�Q@�"]-΄zҊ��S�D�3Nw� �+:P�$��N���9i=�iʅZ>ظ@�e�1�������zB9��^AX���cm|U��7q�'������]L�=�;3�p�hyT��H���	r��A��jȠ��#uFQwQG=�eV�8�0p{D�f3������l-�ETt�w9wZ�N�ݍ9t}R��L2�Nr�Udʬ^9w�wK����:`�,�����8�&nBù$dY+{�+T�����"����jv�c�8��Ԑ�A:u,s	��gT��7��4�J��S	ea���O�7��9�%H����๏z��NOյ�|�ʗ냲��Q��o�!��'�w�o�ߏ���G��}#���,���@u��e��1�c���7�~P�r����y6CQ+B�-g���.XQ<{~��wv���G��)o�@�F ő�[p��|����Ē6?
 v��S�[�R�=����T�T�תV7�^*�)�z��ׅ�D���g�COWǉ孰d�V����P��2�R�$�$^f���0���(#]n����>��ͯ|���[8���g����P�4��v]9������$�D0.��G��;����2�~$�c��*~�Û[��8"?*�0J�)�/XDYն1
gS	��#>��]7|�W"_4L�Co�����.�-��C���a�S3\��4#R�L�Y1�����X�<Ki��q��e�<Έ�ʁ�UsE��p������㤜Ġ����up[Ǳ����B�)H��х��o��٥Z��~d3`��E�;�p܄���G�|=���6��L~]�C���h�4��-F8�K�卒�Р�8z�U�6Ђ��&й��ZLNp���\��ZE�f�~�1��kb�,9>�)��_�*��\Xd�;�K��x_]X<��.[Y�J	���ۧ桟����U����C_"�4��X`�
A
a�;�ƽ^�V�r$9�m7���N3Ԏ�&���>�_F��iQ
�"���U[>�iɊ\��X���G�k��5�0�p*�v�w�����U�9�KJ=�œR?{#+�&��`�ְ}L�J?��K��~'�68 	%��<�ݘoC��.[�c�A|m��e�k����H�Zx�}C��g�se��k6Vi�¥\����\W��%��'���<<K�u-�جzBpo��C,�(�;�����pV�1ǳ������|�}#:��Ú�J�_pg��`$v�Zr���ϰ���!lc�>�uk��sA���4Af�T��xj]�w�CM?!#��aՂ�_�^�R�d|�L���r�a!m�W����Gt�c����1R����Jc�+J(�=Ԏfl�*���]�o����Q�%[~�.yg6J�Q޾Y�b�������Y,�jXZp��)Bͩ��;�����"�0�ŝ�����؇_N&��R��W��O���3�ۑ������]���g
�_�J��"�yd�+=F�.B��%-�J뒬|�+��>��6�`s�����ܯ�3Cb�����$�Pox�̒sǝ��N���#,J7�rzy�ሗ�+A��NqЊl8���ƀ��/����I<9���E�n;� �{[x�0�_���ҝ��1�r��AC���w�L4�|�I���D�Cq������z�,�s��"���Wg:�a"R���Ң':����l��J��D�0�`X1+m�&��^�Q_��0xA�<Xuq5�<�6�|��Ε���}8�,��y�=�]5Wk-8�fs��z�y�|���)��q)��Q���n��aף����M��؋^f���o|��X2��y����x�I&��,TH�i7
σ�i�4!A���Jգ��4��fa���O�\w�űS-�jH�|�)^xL�Ǹ\r_͖	'i;�*M�g��jK�sn �ϔ@�'.5�N�ELc��!��uX=��ў��`?m��^�f���ގ�TM|�hUmQn]?�����3�PD�Q�u)
c.�K@�ՋS.����ω��6�HTz���Їx�1	%ѷjČ�F��S�k�����9õܘ������zw`�K��R.��0���?��Q�)��<���/��q�M�~������q���TQ+�ll:Y��|j'�S�z?�������=</Շ���Y��PY�E�a������z���$��@�G��~uUH�6�YQvn��JL�Єm��&�[+9%��1\t�7j{�?¡�R�ve=���g$F�L}����r�Τ�v	�����,q�D8cU_L�g�$��z��	���P1�����Q��,��t�z�9��0��d/�<�9�����^�77LDV�K�el\Uhn���s�3f(ƥ��;�q�\��o\k��j��@OB��5j3�����Kk}eO�� �!\�� #�wn�$���0���P�`ٞ�@#�^� ��-�tR��v���� �?�*�t�4�y����q6�s����4�p8}7����,��>t�Kl�FPY��_v9��W8�I�&Q#~�����ͼcM��]���_;��6ol�0g~��̾�7*����.��o��.NN��)�0e��3��HV��^�1 A�4��񁖇�����I6�=�ƍ����<5��N`�5e�.O�����S;���_Zys��_Q�#ũ	�e�C2��2��Z���Y��Sܹ1h�2�am?eq%jU$^ FtU���7����u+�3����,`Q����W�a%84���uo��"��ה�c��k2AQj���/�zHk�5M`�B���8�*�Vh�`���lq��Ryj����*�������W��i5)��*6OIɳ�^��ߐ1�NR��[� ƿ¼#�Vw0�m��7��]Z_��tOb�F��ƻ�����?Cr���ɗ�5aQI�E�����>Ѽ����	��E=""�H���S���.��Z��%����{��tT� �����F�9^��8}z���U�L7�PL���3�ٱ�jlM_;w"��С���ᰰq��C���F��+���>;��;����,����	����87��~G�W��Ф���ɨ!�|R�� `��7ȩ�m��8q�`P��Vڧ�n̍�`��b�
�)��"�e�n��� ��W���[������(;��R�>��ij�UH,l�Д�QN�PPcH%���T	��Z���o��յ���K/X�fk�/1.Q��k_QG��F��Z���Ӕ��1Ȳ�^��+�_�fq�&(� f�Y���fM�;�zVQ��)m��uP��M�ʇ3N��a�Rˬ�n�k�|S�z],ǖr �G��K��w��e�����G��C֑u��K3�)���>n��l%M-�n��\�/��	ʥ. �=�#(�#6Łja)���`e|:�n"T��D����y��b����p�q��d�+��v�D��b!b�8뾕�s��j�^���f`�v��vr���Vh2?��6����BՓ�{���绁
&��o�z�d'�"d�N��Q�D���p�\��o.���iy���8>��8����g/c�*�1��`��;/*�*�>9�J����u�U[5��̓i� gy"O�g�5p�#e_����T���++�g���Ƽ���_��hy��@���ʅ}�>����硻F��ߌD��p�6DkxCI(i0W ��ۀ>A��P�fz��l�z�?�(3 V�(ot�4=�{�k�T����$���!���(*�M����c���|�S\j�z�_�G^�g�
 N
HT��=L�"j)�ھ���Ĕ�}�t
��1�E�n-��o����w?�&�X�i<����LJ\����\UN�W�kʰ�C7{ׇ�u��J� g)]���#�|)��')���m���E�;�b�M�o��}�y9�Tc�a`F*��O؝!�*����t�R7�@�d{�W�r�Oy���(�IZbD9`��<�i�����+���L#�wUkk�QF��=7�q�G�u^ׄ�-�	֠�P�B�ɠk����bb���2Oj�b�w7��{�={��Y�]��J���?G�jp�������^7�{�����Y��A>�`o���9y�M��@��-��^����-�o�w�u�WL������3a�(��+��F`=�ǧ���]8���U�J�3X��_�@V�8Mo�&�� "�t��`C)�L*��'�	��B������vB�I��%�*t�9W����a���t��F�;煼 �`t������o�ȸ].:Ѵ����êY�*}���7���^=����6D�WCB�Ԛ�i��,�w��f	T�J	�u��������?�o���l�_SF�z��[����D8� ��}��~B/��xgwk��&7�k8�v텾If�f�ys�9����ג��I�������E�K����z��X�au���W�0��Ę'=��j�.�c��^�M�H���(��t������z�¤�}里5��  �bN�9�F5�T�F0s-�.�s���!�7uYf��d��W�O�������_u5�)F{d��5#�����=�˼�t�+���q-�-X�Z�cF�I� y黿�d���+�E*a3&Xgfl@�gr����0��Fc�6$�g�ni������#�+aS��q�)�R�\V�<䏎�F��گFk�0x�Ȣ劥���1.��le��\Q�����Ln&?i��^ApD��w�x�����ѾN�?�w��
��˜g��v�����WFT@0�cS\C�O*%�Tۣ�B��c�d�U�g!�!]����ʻ�)*���7�d���\���YM0J�S��V�u�l5��!�:ԡ��~�5{��7O��'����z���M��ئ�]y��.�2��(xgk���0�E�jPF�SUE�
���ol\WM@�\�E�����)�������S���)�F.G�۶��~nt��H{��͓�}� ��h �ʥ6��}�2���lv]�O�>S�y�ԭ��I^�|f�+��Ch6��=�£�9��O��8?����غ����>�l�f;g9Q8Eˍ��J�bP�o`�d[��å��aa���1�.�U^ż��$1Ѵv��
Deu/���\7f�29�w#�R�.�����D�H��`��3v��L�Mx8������>N�.�:��+z�&�{w��6�w��������_lD����$d� B��!ƈ��YO߽�r��m4�������;�Ҕ�[c
?:����3�J�������T����lT-)z���>�YYV�)�	F�O��Q��!��W�.������.ڲ����e���\vF�U�jl���s�h+���|}���e��Mo|tkꋑ���$Ѩsa�;�
b&e%M�U��h�<��#�(H���(�ܶ=̿L,����}Ų-
���8���UPh���ũW+���.��ٕ�P8�a$�v��b*Pp�BHv�o�8��^t����15c;4��-J��M�NY}n��YP	/ܜ1P�,a@�{����s,���\�r%h癘%�#�oe��9I7��t�e�H@kw�T�Bq�F���w�(��ڧΡ�r�p�!Rӵ�D
IA3.6󼝯����jv�D���ۨ��bEŵ&�PQ�Hݭ�Lm.z���j���l&9���Q��0�ZY��7]Gþ#� ]-s[+����U�N؃@Y�5���_;'�"�B%�/�R��-4;����s�����\��4�l��	�^y�5S�����)��8����?r��Rً!���=���ܻ�����@� A=����n7��3��{x����=��x�!��E_�G�Tqb�0����KF����®�lM�2�f�͸�
�ns�+�lo�#RȭqhzC.E��Q���V�q�<��r�#�L/<"v��ܘ��o��i��E�CB�{�2 �005qY4˳X��^L-ާM0�ڠ�_8{������(��{	ԲB.������њ�?�rn.^��2��MfZ!1y�->�P;w�2i��
��MN��� ������ZaM]�� @z���ԗT���dETQ�ѐ|����ɓæo��D���y-��ͅ��7�`c8��N��y�z�-+���i}����3\p���_/dQ�a�R�N��M��O�����?�i�=�';8B\W�zqJ���J����=�aJ!���<9�<c߲�iUx]����+6��b��4K#v�a�j�Sxo
G���oc��Hi��d8��~���-aW�N7<�ml��|>�^�����p�s�(���yA+ki�xS�k*������*��3��/~U�(/�KEFf�Ş�⥈�J;��7��q�)����"�E%ȋ4���ꨯ2��L�1�����zzOe�0�=����=AP�[O�᱘�c#	��h�麥Tlo��R����O�P�  &	�Riϻ�0���@[s�B��X
�Z˷n�j�22řm<� �va�������_�~
pt�J�#!�'���%�)��2�NV!b<Ж��J��C�f�@�g|Y�-��|~�X۵M�l;��˜t���-�9���F���8y��ikŽo�6j�y�|JӋ�C���ϠLH����zy���YTd�97�)�~ ���e�S��+�0o�T���t� Vzw|40�MC����d{)���YWu˭x`�b�g�!RYڻ���ַ:Ѩ�|�����@;qn�zh]%u������4�˫�1��8�HO�QI�T���zZ���"��5u�w~�SbxHA��	,U���&t�Ja	�$2�j;�͓���3���=l������)fw�C�q��J|���� U�1N1H7Y�u@n�X��H9�PH�Uj���̞}G�)�K��M�1��,#��� �!��Jʐ0���o�.�<�Iﴮ�gq�i�0�:�����ʓc���o�~��p:�]8P������,¶Cz�=������u��^�+ɿ�@�o�,��L�O�ǏQ��"U�MC����=����8��^0^�e����q�T��,"(��1��^�
+�s�0;�BY8'S�6u�_� vou�����I����O:ҟ�O�KШ���ͳ��`Q��C��ݱ�B���(}	�v����ק"ނa�~RU$K��ڵ�[�Da1#K՝1��@��)�R2�4�w��{����B�U�<�;��1�ؚr�p�S�܄	����HEl��6�3���ˍDS��i^
d�u��%n���u�41%� �eO�W7��h�m45
l��|��wa���s�t�*Ż���QV���ݯМL�����%+����1�B��龍�{W�{����0#-D#.(�M����gi�紓
5|y��ph�a��fXݗ���|�үM2NN���7M�##�WBJ�_x?qDsЙt_'�C�, x4B�T-y���3z�<g�K���Ù�u
���L}���d�Y������h�.\l�ת��L:?�d?݇�3y�THqo!��٬.+۠,�c��d�lJu����2��$,ҭ���E���t�	�B��V����
��X�/q�����*��э�Qx  }�i��]�.�/���?Ͼ[+��BY��8HK�?��Y*�`;���ж�&��7ܪ�hw�
cq��ɡ��0�Q�?+��"���K >��E������8�����<�8sV���g��[[	�4�=1�7���X���c�j�_��L�6Tc�����dR����ȎC�>���G�(_�O��J�66|�<�Ad�n��c �M���m��K7>�H��z��p�X��c���4c�d������u~w����TO�Fs�YTT��Z4�%\�+�(��|ް��c5�G��hM0}�4N�~U����]�d��=)�W�!��\�r�ŕ��rpez
s�6������#�K�Q�&��DB�r#Y����k
W��ߖ�h�wt�AZ"w�n�m�s��b$g���TW_�������f��0
���!D"6�Q�W�I�b�)�oJ��ʙ�
��5�2��-&�3B:f]�%�y���<_��ٻF�;�¯�2d�o	�jѴ�����j�T��ޮ�0ލ@��������S6�$�[I�k���N|�,f��1�Zd>��<���?�&˖!Ӷ�~bH��uI��kՊ.m�/�<���_��R�/�4�a��3�r%:Ĳ>Ѱy�[F[�1��17��í]rZ�V�4��}�m�de��ěywO02�o��!%���vU��;��"���?�j��`��b�OL1�F�T��t����1o�{H�KI���o��;��X��"l	� �"n}♮J=C�㯉�?�\, ��=�W��B/3(82%��3jT�վnU�W�ї:�JI�;��dWD�|lQ6�&�衠��`�F�:�L�v�`u��'�P2����0���{�RF��"��7���GIR��v����q�*	qO��6�A�˗�k*�$i����2T���j��8mL/�����l���R�:/�G"��qC=z�w�9��UrGf���W�q9B1p�Iz+hS�N��tna���pߐ-A�0{� *�P)F/-��S�6HVm��OC��S̭�`n٣訿s.���U^��$�h��3ͳM.�$)��^"n�h��ڭՔ-������Ϧi]/�Ą�m���_?����H.w�����wwr8�lE���iRrߙ48�����z��r�7�<П�+!P�g�0$$�9' �j���gosF��"&�y8���O��/�=���U�hii�
���e', ����f����^$��#��S�61[C��f�� �p�s 	o$G�W�����<&�!�Ke�X�(��z*j��f��ES���J�wU��s\$ UN��|��6�{;/M���y}"����\q���I]ݛ��e���p���ٽ3=_h�9pJ�jCqoy���������R��
�Uq��ϛy�Г��S��R2�vr0������6t�@r@�n�U�[��R�ˏe٤�,�Mߴ������H8S��[�z��������c,�"ᆵ>�y	��5��h���6'cg2��$���^��/s�z���\�������xy�E��:y`�cç�a����(߁ �U����)>��g���W�C\e�񂠨��d�HxtZո�� ښk(��g�CR��Z�ɿ�k��V,�vP���A��rrS�e�����k� ��p��Cʮ�y���I������S8	I��ESu˞'1�Tu����=���hc��[�Ϸ��Z�?U��H.v�����
�pЮ0�*Ne3��<!<Y��J�$���n~�N�R�4r	r�ń��Y��O�U?L'�D��Y���,ib���y$����f�X���H�S !����E�(���H~�s�t����2�-K�V�a�IɌ��߾O|�aez�|��V{͘��xW6�!���:��՟�[���Qѭ�r�~�k |N2?�u�JOH��I�(~;N:��Pڽ3qq�˕���_�Ol��&�D#ҰC>��Xs�����l0Q)(��j��R ����0���!�ƿNέT=�l�'�e��/��+'<M��#��8x�\^�����=ߍ�*i�$@e@�Mk����/�:�Fq>�i�uT���{���2��GC�Y�0�N��9��^w���[c��m�$ZO�.�N� ��ߔ�1�!�%�w�B�|zЇ7�6"}sʙo{t��B�0�-D	�mY=��iep6�H�Q�o�U��<<���~�������jd$�H��vO��Ë`�{�LJ�q� ���"��ܭ��44n�4�?n�eY;_���X�x*yJ���~J����!�
謒믏��0@$K��%��ڧT�I.�?B��*�JC��,?|yw�������vjy��h�O�-�:6Y�~i��o��	�q#�o^� %掗p��y^#�39�8����*��|)q����2����hY
���2R���J��)
��c�v��jH'�(<8i���2?�$��)�0#u���5����^�\����\�D��M=�O��b �fuMEK���_��:��v=U�e�[<�8#(VɈ�1g�gL.���"�����>�2q�ϳ���i����写�#���]�FH0;�`5t>w���-M#� JB&ڜ��Ǵ.0���|4`�����zY�,t5�CI��SU ��4�T;L���P�bHo�m�%u��H�]t�T���\E�oi�c
Ww8QohVU�.�X��E���hb���8ޜH��I���o�!�:�hK'�[ (l�(��}����&cr�f���Ո��3�5�z��b)�P�������G_������_VY����㕺q� �_k��N�dd����Pa�%4v�٦(�A�ۥ�T����A������G~;䡊J�Ӝ?�o�G�ɉ�aʄ ��6,�o����DE(�S{g�]!�I�X}���S9�ܩu��t�~rU�6� �e�Y�"ǒ��ީ/y����YuKi������Ȯw�t����4����A���!�������W�����|:�{l�?r�e�ګ��1� {�i� ��`���@�;�� �0����:���4��(C%��-����|����?�
�c@�#�x(Ϡ>�i�Dj��Ű  ܲ�P��%���/�H9�3�2Q���p��á�uMIѠ�d�b��
�z'����D7��+�#��o([G�S�l�� ������Z7L��1|�j_S�xY���z�*�E��-��C���tV�&���@p���R�"�7݂ ��,Nm�1���ً��Ա"3��,�v�F�P��O�����cYvH�u����_4�?:��Xz��.u�@���0r�%���+|	 ��1�������<
���
�b�#�<T�c �;�Y-�d<�ݓ��~�)�R�T��?�>i�3�0s��2��q�A�?�EW�n5�`��6�cdY�BM�%��v��6�O�,�X��$'CEO�-!�@8xA�2������Z=GM*���9�Hȱ�nHp���UR�س�w�L��r�k�P���*B�G+�g2�:ε7�:/]%LU��W�Q�"mIo�Z�ݨ�l��s��C*)��1"���H���0����.wu�/�z�͸����9�I7�-v�����{U'����q�_�y ���M�/����Ǜ��q�^ZK�6���bɨB��3oN��r��`/+������pܟ��:`�L�F�}�=�*�$)v�h�& 8f��
�f���sk��E�y��[fb5]6��g�|<�t�%��Z��*c[�@��*'2�y^9P	j�H|^(x����ؖM��tSΥ�1�{�F�%};��)��Tkۘ�H���6(�9�-50u8�G����	;|����>&H��mXۀ<�U�n�����M��1l=����Z9�ڷ�}�:z#�1T�:�t1��8���i���a����I�WZ�o��A���}�xe��ѡ,��Ѯ�8��LO�EU��vj��V��$ǲ|0@����jO��B��MX�Ao�N.��N]�jV�@�����fY������8�e~�/\1�]������4��w@ֻ�ʯ���e����>���&�Dx"����܅.dDKC�RL]����[(Ŀ��aߪ��E�۷��v�@N���P�$I
s*	U���_�"�I�n�0��V� �IF���uM.R�Lkl;\����1[�R`o�	bm6��:q��ž�w[NΆNw����)�}�$�Q|�*=�M�@�ʃ���C� �W�D�^Km��6 ��maUM`5�����j�tD�u�0�+}��訵�*߿^ �Z�{|7�%��m���j�z��>Ɲ��c��!d�;mI�9�RF� CC"Φ�/9����׈A��໺M��0�o�NF�M q��ߋ�Z�-��#њK:��\��+[0�ɼ\0���t��c��*��ȯ#9�5f\���>�o�%�@(�' ϖ	���N|C0��Pi~ �kD��U&C·Ɵ�O��PE�|~$�����C����~����㴰c�&Il��ZH�a�/G����G����@�������OHJ�����y�Ti�,]�%�m�t�/�����t�xmж�.I�)D��R�X+�X;+;hH`��|%�7[���+}��8�M�#�������:�)��jG:�����q�Fk����Sڢ8�׎�4O�z��V���`��mY/�_9 �x|4]&_���������f��B$������/^�:G�C��Đ�AGl��Ǧ���=�����Ƥ -4WCx9���5�&1�w�(�&�n>��c]�=Y� ������*�?�!]��&}c����x�yuEdV.��:�s�|Y=�o;c}���<e/�=\C�(p5~(��I>Ѿ������h���!7�X��m)яr���Sk4#��*%]r�䄬V��Ã��K������T�Lݽ��N��������ۊ���\=��_T�����@��B>߻���YNf��*��!��B!�`��n��IAc�k#u'!���Фab���#ju��$ ���x*��?BXB�8fz�������M?:���5Iڊ��Ǎl�³�n����0�¯6�((�q�A1Ú��%�U6*�2�# �~Q�02����Ӽ ��xR�J�M���ae��yl��w�fz�M��o��j�Q���-=k�3!=:��rM3C$&�B������q�	n��u~�ey��f���r��`u�wfS9��l+Ľ���9�y4O:�'*N���kRO����&=q[-��0�o�Y���De�)Á�>��2`Ij�w�^X��;�>��ȌM��mB��bE# �r勉��G%5����P�!
}�mR�E�h4U�N�����h,��g,\IvQ�N1'�R�
���j���ŅF!���@�V2X�ăHij�BG��*��d�9�5.��2�L��e�I ��KJ9v�����+��P�f��&����CF(��=C�lx?�ᒳD1\�k���`cID=�[������b��?0˦���=�c������W6�,A���SL�yC-�I����d�;;����[�&g�3}}�$5�7�I2l�z����|ZǢ`v�23r�e���M��Î}�Jf���FJ9���Ȥ|p�w8q�%���a�8����܂d]F��V�V��뱜��V	�p�̆ķ4,-��-����p���h��eFF^%/�� �f��us��%x�8�c.6]�ȗ&��Q|��Be�-�t�M�>ҕ #��
�+4�r�
X&�Ce��/��/�sBđއ���1��d�`�N����p��� E�Ln_	��M�&&t�zk�2�Q߱u�8�V�W���Xe_U����8��D���`떓ݨO��pP&V}ؙ��K�&�?k:�{ZA�M�Wݳ���df�����W�#i�6�&�Yg���L
u͙��6�w�]`����c�$&OY�p:h��E����2��e6��[��I��.����Uj��2'�A����ŭWµ<���Gm�R�|ngd�*Z2�ȸ
��� ;�9�	���!�>B���r�&h���v��+���X�E1_B�<M��n.px��x7��>?Ћ:��&���"V�~Q�IeC?e�K/��y���̢�<\�g������y�oV��7�a�+rN�~���n$W�'��ћXH�~� 
d���BO\�=<dΡ.�TE���ֺ��|�KRÒǱ'_�i�����!�B���PFG�8*�����Z�+��T���N��� k�֪T��f��n�j�%/�A��o���s���|A��u���F�*z�����(O,f�� 怒��?��k�l�/X\aƕ^�j2�|��4�N���|G�h�z�I/�n�^ja$��Ly���:"�sQq�H��g�[o���/k�=p�W%���,]�s�Tfl��(���x�ΰ�GѐoMKG�\��1P�6x��0ox���[7ᆵ��g�����T5�>4X���\��A�./���.���Zk{��J��57�߂�� ���]h*T�#���ㆽm��xnHh$�����^請@5�*ˌ��������n�#�>�e�9�J"��% ZrZ�e�J���vL��Ɉ��� ��L�TqKs��L�.%������a�VD�S}|�(���0VT��y~�PF*>A�e�
�.��)�v��l*�re��^xys�����}�c]<EQ�e�X��P��"���!�������GZ
�33}m���k�UdxaT���r�:lq����o�:�TDu�*��,�"�jnq.x�{�8��)e�bK�d
�k�HpW�/��g(�s�H��}�CG�ytE�c�ѻy�����C<��+i�3i<�a��|d����lxW1�ӥEU޿��a�/N2��tG'�r�!��b�Sh�-���^8�hȇxT��T4��gd�P=w�����?�zo�Ƈ'!�ku�m��t�;��v�t���l}D��ǰ�0�gi�kN`���ћ7g�ۋL_~�5��e?h��-��+�C<(�<'v���8���RCc�x����y�����))��dO��Uc%�PEm�}[�2�V�Cn!?�.�j���E�M���b��(��'g�_WX�1{5J���"/�6��k.ktWI0xQ�~Q��ܮ�ǸpY,��:�+TJ[�>�LP�k7ud�����uG���ju�|	�����/ߟ=$ḷ�`#��^�	�BH�6EVa@��(��W���/����)�Q,��WZ�E��MU��� 
ԲL�u�!������h����-ذf���$��T�B����e�����.��pX��ߡ�x \���X,�]�?�\��E^�A�I�f�;��e���Օ��C���4����}����G<j��G�ŋX�䄌<̐p%�k�4c.��/H
F�d�'��$��3����(��x:���[� �t^�k�	��mUͨ����X�C*>�;R!�o�%��id���[m9�S��8VwH�#Ů����:>�µ����ŐE�U��y��<T4+?�z���ӽ��ci����%[SŔ(hv�A�P0��L�X�-�6=�3����X��� mQe�ش�ʏ-K��|�����X>ɻ�붅�$�fЩ�M�:�U��#��j�ʴ�o��HwG+�k�(��L������Ki��qB\@5��Vp���yRW�����}"��:�C����� B���_i-���x�xB�����QT*��㋃�.J����)b��\��K��75=՗�����4M)�x�(�(#�C�5^�O$O��X���B��g���O	Q��r^�Nϳ�ir� :0���HI��Z�f��hl?<^)vS��?��彉Ny���5��5!@�XsDdT�'�L��͜��/0�n"�;
\-�E��x��~�Wo���gF�	��L���Og�[����O4�ٷ��I��f�g_��%����U� AeLv{������ e�'��`|�QH��v����h���Yq� �Ba��xX�����g��mr��$e&�*��с�3��(�kv�*O�?�0�	Y�����{��1c �c�te:�0���ɒY���e����-`�����L�a�[\�;g��Cމ�%�tσgI�[؍9��J����ֽiO&�OV�Հ� �P�C�Z�ܫ�$�-ԥ���D�e+�*b+�R(8��	�v���9�uk��$�[�EB������ng9���2� ��۞���2�*>T�T�����:<ƙϝ����~���[8'�@�{O¼:�rHv��.Z�e92D!�=���/�;	-y.��굻N�<�f4LᅗAk�I}�#���{��[W�1�@!��H�[WfiF0@{0���ͤ�����8Pm��ԫ��I�Z���n��a.WH�a�� �vt��W�k�y%�s�m��4�b�(����n�"������L�"u��>M���3�)l���a�@O��+�:�t����<�$�:�Ŀ�Xf=p@�JaL3�N���hg�Gu���z�x�
D���!�tzB3���*�)��|`��*��<��e^25.���~����r�B�K��k�Q�7,������F"3� ��m��=U��t�Q��� ��d��U[�L�v��3Z��嫶�:�Ki�ތ��6�
n��z]��P��PI��R�0������W�օZ���!*���Q:6��-�\��+P��st�l��/і�����6���ъ���/F��U��;�,/Q��n*���,��+��c���{U��m��~I�s)B���w �b���Z���
���h4pu6a7o~�"��O:5�zQol�F��,��& Y*QJu�o� �^��U,<4b ���-�O�H�9d�����3�;����.�[���?���c�
�Hzs�7�~M���)xW�H�G�[��Xh��(�9���]Q�v;���C�����<�א$�v>,$W��	�W���(Ya�{&6å:󫉄a���ړ����>Wʐ��!�#Y!v�W7l�L\�1��X��:x�q��;f��#u�T�_����]��~c:Z��:!��+H����ǲ皡(׌R	h
���^$2FjHD�8�I�OuHB�L�����h��_!@�(�t"�e*��ޔ�lu���2d��$�s�NxM�G��n��0G����]7b�\(�oPZ�Ne|�8�a_��v��3���R܁E��_���F�Sy��X7�No?D4��Ma����/j�í�6��1w������b�,G�J��4<�����y��h�S���~g��Ƃ��
�i���-���)�[=ν���c;RQ*�]���IaQW�SH.�����l����*�-�0���*�g�/��%�VQ�ڡ��2�3��$�]	�`���q"²D����r\�<�Q��5�>���1d��2s?)�Z�U��d&Aעv��=
��� ��C?B�?(�'��S�f��H�H���=�FP$�����M����]�15��-��UJw6��:jL��z���$+�շ^~kh*Cw�@�^|�(R���M��Bm,挓�=�;��Ȝ(>�?/��P���f6�褑%�k�����h_xX΢��}�)���%�݇fP�[Z�n�0̝Uۜ��ys�S׳j��&�&}M�����b^��3��������@��_���"� O����~`�)���|��^���`C��������҃?��/���4�����}��X��7kl�e\ᾉ�=��$�P?�j��FP��+_I @.�r�>3�c�[��6û�))̹��Pw�T��m���|�E����Y����|�α-ɢR���d�e2���S��8����8��(��g�P����&g�3;�Sq�z;�^�eG8)l��j�J�bbs�}�P��1Qz�y�B��Ԛ���f�vZL�qe��+��N��:�������}��Ө�Te����P6�נ���nM���h�E��|#�Z�0�wC�M��'����[3�*(��7+��Ȏ�`�^��Oai����
�t@2��LB��.H�r�u;o�.���Ǵ𕽰\>NC�`ݶ�3P���6䭾�a����7���Ҫ����Ї��"Y 	�9́Ȣ`��܍y�R�~���evV���.���ZS�$ݏx��%�*ò*��V�LQ��H��K<u�\�
�U]v���z$����?'_{�"��k뵕Wq�
�!�ǉ���P,t獧�C�^��Ъ}�+%|�5�L(C�b��@�D!}��o�W|RO�l!{������ �n��_b0�;A�6r	Tܗ�Z:�z�q����߸�����)�!a�Ԗ �qұY����s���VO:oel�'��Y��2����T����\]>6��/��o�nV��������ZX�~����]&Ƚ���5�	��Q��V��1��_Bŉ̨�,�v]�˽�}��C���D����,U���=��5Xw�1RA�7���	
�c/G@���h�������05��:�������*<d�����	���6�F��'s��/>�҆ݣ�^�!a j�_�WD�ݍ��9=�u`�� ���si-�����wi�q"��#"9��1sV�ߝ8'_K>9X!Oqr"���.�"%0>�F��9(Q~:@��@�&2閨�����7���A`���c�;9�I%��[g�q�a4h/[0�ҞU��=W� DK޾f/㹔ʷ��HNOӸŴ!h'?Bf'�%gۂT'�}�<D���Fa�T���� J���J��QP��W���E0�B{�`��펟���Ж�'t �oK8�� ��9|��0�0�t\��k�?[8�_�s����9��$fLn���h�b�����Y����Mtʈ�K�y⢅@]��$��!�@i��<�P	3�PΑ�6�Es���>5�F�ȃ���r!���[J�^� W?����>9Ïl?���^�fآ�����0��<yI���t�M�N>�ވ�k����y�r�J{��ģ*+r���͇�*<>�/+���69.��o?4�>H�+���q��	a�l� ���X���Q\��)]��9�'/�1[�9p^���-��:���׳�ׯ�2�O{3�%�4�n��"��y��qȉ<y"�H]ۮpqc�.R	\}q`�u�����Ψ��;>�kN���7���)V�2;��I�4y�R��w ��;�a3�]���ۙ�}�4d�T��d"����9��,麭B�3(�Z��Z��b��^_�����+�8��H� ���p�mfl��U�h� h}��(���G�;����Z�1N6����9�i�!8�3�)z�%D���a��� �;�����6�J�J�j����HZ�چ��ă���т��x[���W�UtęǇ:~j�qAb�X`ž5�*v���������5d)���:Kx����i�@m����/�	l���J����a�6���jt�R����Fρ.M�c��+-*�,&D�l9�Cg�*��I���ȝ�I�L?��}��� �Mo�P�Aq�^�����Q$�����뤯�)X����Y ��;���������-�����|R��5^Ul
����Yg����pZr�hм�|�,����jh+N`MV5սA,�8�&iW5�P?;	���mw��p���XhUC�TpN����h$�׿�&e�Z��p˾k:�����0&�T�T4n8���&&t�J����v��>${r�(�u�!C#Ҏ����,��Ju���@�� �� �I�y_��%���r7E9?>T񪜻R���ܟL������OtY� �m�"}�ȧHbZ�5���ϯi��	����Q�L�Ϊ�S�NR���}�`2�ٽ��֤�J����Q5��y$��(%r4�4q�.N5�����]��o�/;	8ɢ�&|XN-s(����KxO����u};����{Bx%�
t�u̬ ��ռ����a\=4�sy����U�+�<<��������x��
��� ,�G&�i�a*k�F���z.H�)ɷ^��;�r�~&�UVd�ں�_���S��&ӭ4U�~�=L�X�u\��%�\R��r�֤�>)��	K�����A�ejCC�C�����5�i��֐y��A�b[lk< b�><�G�Q��Q�+w��j$��-��/h��XmI
���~��c]���p��H��/fʍ4�\k��k�>*3�x�����ww���N��պ���ܺ��εO�fYSCC"��5����4`&��馞qf��aQn�h'�;����pJR�Kk�e0CI��Ξ�
��#�7�}��
X<��E$��CA�Yg��F�^_I��*�ИaH�b&-,\�N"J�/U����h���-�,I �%�`����\Y���o��J{�	y�,�$� ��Vr����	�dv�߷) ^��G���!�A�|��87hӝs�"T3�p�3���a��gC��<�X&i�6��L=����_���3�G����R]΃	��Mܹ�w!�s��W����.�������Z)�W�BNp��,�4
�;`���y'�)��\���Fy,=��v='JN��o��#���
��
i+�^&	a���B..�($�РW�nJ��r�tRe<�d���u�]�1��z)Lc;�OG���7���J��Z����D{-/��o�Њf���,3�
GD� w�qw&Rۦ���y��ܿH�q�0@��O̍IG�H�)*p�T^kRM�h/�Зv!��"��T� �M��E��K�,���g6L��pd�hX ���G�P��i�ꬩ���<�L�d�mS�����@VR�JN~ � ���	�I��I2�2>�=��=Y�_��#�o�O�u��i�Y1y1���R���g1�f�3���9'JF�r&�[R���qEv��b�L!���ȃf���]Y='�����e���M$߱�����t*:�s>;=��k�?�,�v�ש#�9��ӧ!��Y���
;f?��ǾDF����E}\���d7`�{B�(�p�J��E!�ƞiG3�t�������+���jѦ~j�c��$�~�W���#~m��+�>ƕ�mQ���7m��}���+���	j=>��Qp����|1p�S����O���v�rf�A��ķ�%u�WN��[��j���DӁ�t�>��`�������~9�������DBb?SH<d<���hI�C��O��Ҕ�h�0@�_Z�+�~��G�r hu+�j�!:�Ҹ��Δ��!�g)-/f��s��G�]�>��4�$�Zx���9N\��%�Z�I�2�9�^=�3����� ���M��2���n�趣�y;�x�RN!b����\fy�Ϫ�;�Y���I:��(hyt8�����o>�{t��gq�d&c_ k��Fh�0�l�$���b�?�T���u��=��o��|YF����T�2�[�8�*���b8��>��go=X
(�聾k�V�7���C�Bcd��~*���#5�����̳Cq����/�z��h'�bWf�䐝�&����k�����ՖE��z�DB-c�U�k�|�!�9�%�Y�otI�Y���3O�����+�5F�L��)l�1�_��`Y[����5,�"Wߪ�;/H-Yo�C� ��zr��0�ʁ���]��uD� ~�?H1�д�m���]V@�LtGn�i�Ғ+�'��>��Ȗ� 4��k���T��-w�F�z���}5������i��hP_�{'�bLЪ�Ȼ?��jd��ц0 ~ OB�p�(~߅�*e�
\�ѓ��lv������f<�~�)�Oc�fյt�?T���N��5dh�YQ7d<@�M��3Y����E.�U�5�Le�o�4vwJ�L�������2\h=QX\ވ
�)�S R�;�����@�FmI�_X��س;Y!���0�uU���bU��݇ �2�K�疑>U�"�7��H�������Ь۷ݧ��4TMe�3��4��KR5���N#���@8#!f��{E������6� ��9.M���(Un4�4{����=���2�E�dX��PFq��\UpF���4$\7�̣`x��k5I�� �R�^A4�/Un���l�V-
�`ذ=� M+'��ev�����Ro�7|�ug�|��膗M�m�I��J.��u�$��k���lJCc�.c���A`?4)y�Lͷ�=`�]6�M��B�%�v�:^����nO��Ν��|��4&��Ẍ2�4�؃�Z�Vr���2W��{Ṹ���>M������0���������"8ա��p��$h��Nw-j/��a��v ���I�����"���#Ԃ�P��YM��
���LI�L�+�}/ٝ�)��!��3c:φ�t�[�P���i�8(!n@��B�g��Ћ9�N�����]��`��VL���y�0�;|��kmU)Qi
jL�Bc�%S�\#N�F�����q=@[�
�"�������쫌 �\sS~ԗl�Aq�9����b<fP.(����;�����m$>=uB�T���X�e`�%�s� �b����#�r�"+�fUL��-���k�O�C�B�<��2����M��t?�F�ߙ�رYk�+4Q�<u���^M.K��tF6��hJ��#-)FW*|���B����G_��N4��J��\k"qkQ�b�	�����/���l�&6��4�G�� ��Nr�ۓ��<�unT��h�qUA2��46�㈛��wB,��ٓ���$���Թ��d���˂OK,_��O%qY��)xp�/Ԕ���vT�yb�J�߀�_e��6��,����&��S�S���ROqe��AC����pul/?se1�����cⴘ��k�p2 ��J\������~
�Z���2����3V���f?�+ !�2������(��st�w�]��b�ʈ��
Cw��'9�����@s�x����Y��嶐�4�$*�slHi�n�jt�>����Zڴd�!���]�����=�²��APc�/��s���<{Ƶ��T\`�������	�n��+��Q�Ì/}���"���`����
��f4uGe'�u���9��W�L_��Fs�L��aSc&��/� P.�O(f�V��`���ῺF
W�@�yG��\�@-V��0����f";G�E�c��䍗BR�T���=�kt8��l!����/eT����}�{��O������ޤ+��!UqB�c�؃�����*z	}u=Wo$��,��a��[%�aUF�#�@���׮�[�KL����Bk�"�ȶ\�X�}�t�1����%5�_��O�?'�X���g�q�mkA�[��4�>���Ï��!�F�RA;hX�5`���sC���u�
B�!؇��^�H��X���~z��o�\��Ql��C�{eH�s��L��D�`���S����Q.��i�]�b�"�,�#=v�t�͛p�ߴ#�'�Z������%�4v�T|&��$�r8�QK�������y�K9𘓗#�����0�xF��hn�v�!X�`PZ�۳�Y!Rx���mH�>wCP���U>+w��Ƕ}G�'�J;=%���0�}ߕe����@?�G�*�.驣Ä1�%�#��Ce�j�,Y��(u�JJ���m;�l&���`mMy�'\�l��v&�6�2BrMa;aZ0�F�(
.�7��z	���uE�n�9�3�]>�0Fz#DP�k��6%�,�sE4c�ܝ̗LRQ�&�n���t��!��\3�Lr�?P��?�ށ'�§�bK+'�:!�I��2t��s���p�
et�|Nܥ���_Fiޏ��"�W��)�Rg֍�%�nB���{�/���	���>"�Y����yZ�ÈUy��B�'ԩ���c�bȞz��Ѥ��Rs��}Mw��x��	�cb�n�jT��` �KݕU!W�ޏp�u(f�[�����i��5'�������޿�;�%t�qL��I����$�d����J��5Ju��D��~R�x��dYS!t��LP,�����]�������{ ����j�1��qk9���c1���++i�c�F;�e�P��d�6�g�DkY���\�|�O~D7���� �7_�aV�8i���>N�<����Ϭ�I���ل���u����K)y��ei���Ӣ'.ң��|�d�g/^F�36��i�$P~�$�G�杖�f���C?>̇�CG�s��[�������o��	r��FH0���*��d.t��(7��Z�}|����/�Ś4ˎr�o��b)��guhs8������u��w��J�j����M�>�sio�3�/���6[ 1&�S
����]r񂖏�j_d�#� ��c�4_�z���u�
������cڻz��J�P~�����q�3:}]O����7w��yj�-h���B��Z�J�͟�Y���@�c��s&¬S���t͙��I���0ղ��j�#!�y�%�\�o��,����C:���O4��YwZ=�:{�s�S;��fP�Bgm_��cȮ�g��VQ��V��-o��\�z�}���?}>�cxԇ �v~����@O�� ���dd)��-�����F7�(��dK�I�E�xWN*��P푕:ш>�v�|;9L�奻Ohx��<���B<����Mqi�\��Y��sf�*)������gP�0SpWyst�/)���	�.�|�8`�`��_�ӝ��X�m��v��^�(��*�$�eG����2�~o�Q5���dN��z���,~`��kJ���j[��N�r�	t��Ȁ�����3����A��*����H5��\��o苂���;/:��'�����@��*�<d;���ƶ�9�-,��4�gǶ��C~��������}�C�C+em�ڰ9�����c�j;���Cy��V� ��x��R{�ە��<��NGL��ѳ ��G�;#�[�*�xx)Ztu���#^	���k`PUV],���]m�S��L�͹b���^L�Ac�����;H��蕢x��sJ�^��U��b����$��X��a���^ٟ�-���[' ma��4��� ^�!�q�R���lpVmsI�⽪;L�;- u��e&K/b����y��I �6A-d���T�6"����+�gl�46���Gu�&`u�"cf+, �'pmX��qti���B遣�*��Ը��R�M�#HE2��2�����P2�*`��VW~٨�w��K����2�d ������ΊѮ+��m���϶/���R�Y`��< ,��"
3z�g��m�O��1%%�ﮔ;U�P��;���{V^ʆ�`�`����˓Epto�����*���$~�e�>S����?�F�l�T�`k)�	S\f}F2��w~���ʤk�L]5]������C�WH��#�m)��RQ[����9�=[L��=�5Z%N(��]0��������$�M�����0��A��X�Cx�[� ,�dΐ�g�������g<V��y	�M���
bc��[
t7�P���_�[�C�����a�I�-����D�z�;�X����A^�H���d��́d�韐�P>��[��4���u|u�7��9{�<�z�x6	V:@ye�"*x)�P(R֤��ǭC��nƾ#��]z�'Msj����a��4�(��qO[/�E5f��.�s�B��Ծ�b+�$`�n��v�/�[@d�]b;1��I��Ҝ