��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U����*�6T�C��TR�ji����6,?��v�sR�6ϳ�8do�Wq ��jt�<�����.���L��d��A(�1C��S��ˏ�~���Y���E��nh�oj�[���Oc%� �K�b5�\(�CU�Yp�Ze����:��Þڶ��S[�E�+����i����W��w��k� 8����6~I�<��;�2ߦ�?�Q�c2z�$	H��a�fȓVVR�p^[_���J�pX�M�;���y5A����|�H 9�,�'�����u����?Β0b�Ŝ�Nj�I*�y%�y����C
V�l�_?���@��&z���ڔ�-V(��R�q����ȵ5`n����V}=:hD���h`A�@�R	N�ga�EI���Ɇ�0�~�����ht��m�$S���V�c�<��Ӌ+��}ݜ����]��i� �
�I��Ʒ,�_��K��R�0K.�5=2�ydZ�q^��9y�o���/���4$$+�=�C�:Y�s��Oԇ�^|F �@68�-�F�0q��U[��^�����Nr��+,�5N?
��������&�.�z��T�0�I'��a�I����/��#:6�hдH������X�>�V���xR�x�#�X�처�*\�U&�Nu��]"�MX�w�.u�$���]c�+��SI�$����i4�f�`�'ZJ?�=jq�%� 9vO�Gzo�ei�&�^b��k_c���y��Hi�c���;���J�&:쁬�ۅ�24s<fm�����z����D�O���7�9v��

���ʥ���z-�|O��'�$�X����r�ag钐k�Xd�v�
�d��ڦ��&&�l������Ԁ~K`�Vd�1C�2��)$�2r���r:wY�t���@t 5w?F�6��yw�e�>� yCq�%����:SM�������0l]ey!��~{�j�$���N�3��#��"�J���o�{`�"p�Uw�7Lt����������i���5�k����j�i��±�!�z�}K���9�2P{�hMBaL~(���ъ+�]5K-��b�;����QFrI���i�Ż�_2(�=�zzvtmu�z�@���~��LTR�k_�(ǎJd��Z����zO��+��~�*7�����UWmuC-�@��(A�-A쎢�ipД2�:�oP����� �E\��~�eNY���d^��������ik�;?{�t���Nf�����ܡ1jfT��X`��[��~
�Eѓ��'������b�>JR�贎���f����2�(��j`��	ӝ0~��I�)	{��]�rʏ��|�D��DL�4f�Q���3=k�ޝwR��j�pp�
5��3�Y�xcO4F��sܳ�DX�h�K���m��k��]�If�՗�� �1D/6���.���i@�I�r�Ro�44��g���$q`�B�.�����qb��^W�
(�7��S����Ƚ����>��&��������;���럍���X9_� �:ԁ��T'�)k��"���c�"kn./~I/sߝF�
3|ƀS�!j�"%�'�aN3�Vbu�{�wu�D�J�RS�q��������D��C��G���0����g5���:��Bt���a�S��bXB���MN�nX=ZZ�!J^<~Q��/��>U:Sw&C�z�h���-�;~q�(x	-��>� ����iU�>�a�[�������V��j��R�n�/��䈟�H�82Q�;����.�땨�c���rhO�4��S��i� &+��� -[A�~�G���#��,�������e���q��^�-���lo	�㌗�%�8��$1zu�����a�|Rh����������ϔb�Ms��<�6ˆ�������� Z݆�"�h �nk2�wL��w��X��.侷w�%]pXZ�fy� ��5���`�3OM��Qup@ZV�C&Tx��x��!��t&��r'+�8�L�B��t �	��:I]�Sw}7Y�N�0ԳȌBg���ʰY`��/���WW<�Jvĵ�\r�U&=���W��� J�ȕh�ݯ:��_��%�|eWH8ƘP�.o�|�򯋱 i�i��ȶ��27������d}t���|�AE�I�iU0`�{B�� mP�ف;��l\r&�a��;4��-��DC�f'��k���c�Z"쒨�C�e���|���8+���q���aQ!��`K ���Q:�tIH����u��is�o��h��i��<�kr����M��bī�hBj��f�71,�kVs^���>Ԓ�qv�� ����y��	jp.�u�]%C����#����t��R�����X����r(���:躀�k#�3�p1I�n�Q$��[h��V;�:����)���=6P��S��+(�o�� Bk*j�9RY��J���:�*7��׿0�F����n�w\�99�v�OO��#��g�I��-�{ �w��b&�5�"	κ\�MJ'mpA(�	��S�y��~\P;4����4L(�xtQ:��\��{�2����zy�x*.pG?���̓1s�p��a��$'�n���x`�ڷ�d��\�!�����$[�ؒ�3D�@D��X/�����c0L�>pqu�͑����"�|�z)��2�/��K���wGڈ�����%M<���g�e#���a�KK@���i�8���mٯ��V߹�'����zX-J
͌0F�Ĕ�\oWcu*Ɏq�Ml��9�*�q�=�&�ن{����w;�vW���_S��J ��O��_��)1G��B�8 �c(����h�mH��v�0��	�mc��Jͣ�G8�y�8�����3�����RKX�ik=�0퀲;��Z.==�~��jt�I�Y�4��,�0g�������OKxmp(p��W+��ip=<�T�����d!���	�ʅR�̧�ݥ��
(�e��L��xd��)4K�JV+Ei۸�j.ӫ��"�(vt=�D�/1��@���n-i��6ں˲T7���h��3y��=�
+'&��$��C%Ze�c�:{}w��w�0ʠ\k�98�Gs�e]̕�B���CgC ��I��}�a�	"��.l=�|�	`,=j
�����$�E���i�K����������k�웶d��\r�&��$�4�=��W� ���:�4=�����Y�*`���2'<'��&�2�Lo;Rˍ|�tf7%���5Z��ڌgYѲR����Nv�	��?F��6)'�s>�蛾39e4իKڧ��X�ȂtXG��,�Lo�Ez)��y�*�8z�)d�+U��p���G�����
��0e�K��ԹA�]�Ȩ���HY����vw8˃��SL�i�B/�拑����ߒꬦZkߒ������D�'��(��M�+@ֿD��ӻ� �qf� �a����5��aLE���vX/RXp�
�FA\5�n�Ch*��#M��ѧ�j��<�������\}�
�e� �e��Ua_���w�	��tY �2~��Ee�W8���t��v5U�s����U���������í�`�BE��/��/��A���y)wT	�������	i��E-eG<Λ ��)NH�"���<c-���Ȏ��̰ EO#C�!4�{3$:�m�[iM:�p�2��rXm�ܞB�&�`�e�������R&q�$��[��T��`Vw�D��e�����4�~ɎҸ�#٨ē��e�#�!����]��#E�!�r�>���(�ai���V�,�mw�\��c;�����Z.G�����Mu��X�a�ʭ}W��ܣ�3�՝�����Iz�x���|=�ϲ���Ɩ�B�1Reg~0�	S�L3&�~h�g����D��4�Ż�g�a5[�]|m�ԏO"�z��J����q�2lpL�U\u���~�d���;��3��j��(g��5SSSd�/.�ܑ`���k�6�A�
�e$�6�e@�p�����S��:�K�ڭc Ǳ�-��m�l0��dCY�r	���
�Y@��U ��Sn#�m�Ц�������
^S\���H�E.�h��k7ĭp��GY�����"��K��I��1�E��F�(Ʉ�۰�s\#=�|	��;mt���K����*\��[>�;2ȹ�Αo7���T�����vc8$���?�&�S@�͖��X��C��:7�j4B��zƵ%N���y�3z� k]�7ǘd�枂o����?s�2�j�����BA�P�gA:����o]��j�'�G>�o�'IQ	���`�)#2	鱃t�e�"F��祛�!����4�-�]M!TBY+h:+���R[���(3����^ӑ3=���J	�w8B|IJ3Ŵ.	��r��|��ե������_���0�&^=(�\R���w?F��@T�\*?��O����3�;o����ZK��C
�>Ž�[�кF	��,V&�7��l+H�:Z�lԨ�2�U�s~?������O�����29	�3H1?��yq�`����Y�
������%Z!�]m��˒)�P F��O����Ahoq�҈�#�D�7��rXٽ�q���2������=%��>�n�t؀�F��ݿm������0�K;�ѭq��	vz��w�%�,go�C�;`¬˕p4���>��e�N
<>og�܎�MR|��; �
�t��4N�)$�@=�|��)Xf���ܙ�����G���%.��Z����C��9�N��Տǫ��w��F��x�S�^>'+�W�^�=���ݘ�fТ��I ��,s�A"� ���pŊŜ!Z|��0~����V���P�K�'7s�L�7p�.B(a(�+\��V�#øK&2∬z����
�$P�Q�b�����U��
%����O�f�>��v���^;$�,쫐c/�o�/��L��`:��dU��t���=l��������e�������C��1�ih.�$̫pȨ�ڢY3���p <^P�5�vN�H�
Uu��b�Gq��q�IN��9t�c�2�N}�fgƂF��⸟���7�<������'�e�Gb8ePM�z!�1
�VLMo\����PxW<�?�������=�0Sm֔���$f�E���j\�^Z���n��4(����"��v����o6`��p�o��N���r��q��p�Ɔ/gm`!P+9�V����C6���.x����=|��m�>�I0
����E�����6\��,,@�Nz�]n� �Q���A����8���䦊9֙����ش ��뾨��OD�u�8���J׫6�ps(3i��.���)�Ǒ��/@��~g{1s�P�:U�X��a�:m�/$⎍���K�K8C��/G�"k���Y"ۻ�ܸ��	n��j��ǸO�q'g�������S�a�/K��ӀaE�p��v`w�~��F9ė�c��L�g/�8Ƥ@���U��0�R�8<벪�l9����@��J/�7����9)�!�3i>��p��p~������k���K����؋,�$2n�5�u���<¦F*���v��y�� =|���0�<��}�����\��XC�U,�i<�Eޣ����B��A�+���?�,���_3B�Z�U裞�!�I/��������/�~�NziJ���'`�ڽ�!�຋���a]3ճ!�
�,P��%��)Ͻ;ߎG x��2u�7DM�D�Q/�'�y\z�%��YC'��tw_��w�D��2 rU��,����F��X��2���+0%DS_\�������q9�*"k*\��I{���>�Ks9a�.�+�ƽw�R���=�8���{��.<���_L��^����~����L]~&�s���};Q��X��]�|1W��UsG-�q��A)5�5�����
�V����.n�5l�UMZ��?�k���2W� ����=9c�q���ƪ�t�Hu��U��Aw��Gw��[���%�D�Xq�X��Ҿy�����a�t��zw�! ��z�3萡��P�o�p���v�#GEG���fq�ii�2J�WI��P~��1�.Q"�e�;���M���|p��l�ˡ�c9:����.�T&�5y���q!���vA�Q^t9�Z�g�C�X%~=~*kiP����K#Ɓ�mQ�c���[I��fԠ7�67~�s�lg�[���\*���3|D��V�b�9޳Y��<��2��{���t�xB�]{&� Sh.u�ƅ��)�l�
��8y���s!�_p��<F�ƴټ��Q0���#��M$d��]R6(�g� ���d��n�H1��+����V��c�.F�)R��*��踽��[��kOA�bpI�!��aY��%�mgމ�Tq��R��{e�"H����N��@�/�[Ir	�F��e�c��c2 L`P0�g�k�z�m&��C�R���h��k�;���8p�������SY��ݸHݓ�`ܶr@P���c}�\	��~�:��h?�P[޸��B�	*�?ߞ���s�Dڃp!n��\��V����ZE�7�f�N�>匹q���j���LX���vε|i�%�ĉ,�4�CA���k|%����j�d9}�35��1�H
{��}���M��:��rUY!D녪���Le!6���D����҇�ܽ�
k� �w�c���6=��o~p	�w���wؐ�i�s=�x��C�P7��8�aX�}�������CH��8�)�A���v�E�y.�z2��{I�2EY2��R�w5�*�IO�Qy��ݢ�':��z��5�V�:jǧF\d4a��Wc�b�ٟ���� x�A�z7*�٘�q\J��: �}T�դo��P�z��*ߋ�Qd��p�\���}B��� ~щ��7�1�)J9R6��cu_��V�:0w`{��)̓s�\�! M���)���`6�&,lv����+��Yя��y���b0V�x`o ����؎�O�����P)�fz�͝x���Y"X�[4=T2��k�w1!F�J��DϤ7T���mX�0��ʐĪ��Ů��K/��u�����e��=�}]��/1t.�N�o@�lY�L�giY9F����Q��D��w�Lw���S-��u�6�YX��m��;�i�{�����w��Z���$�L������3�3,leG� �J}�ɻX���j sZ�Ow�E�wuq�Τ;���`wZ��$�<0�@��8���Y����堉��9v�o�Z����9�8+�J�zQ�J�ΪA���d̊�̷+v
���T3߀�.�gy��0"�'����]��c�WY�Le����M�I�#g(����ДK�	�� K�;����8�W�`�*vȠ����e]�[e�
?��5�_c�v��q�>LQ��tl��摒rgTP��>T��znD��+�L�q��Aj��`7Lm�{�<g��XX��]�՞9��q4���̵r�����\#���;���^(꺛�91��L|c�g�#���=mKn�i�PK<��L�������C>��Өl��m��ҿpT*��mX�!U���6�Y�,:���=�j��H;̨󩚒�.&͗w�Z��L$�Z��t����@���Y�҈*v���9	�Ih���ܤ�K�7�8�vm!KJ�y�L�/rP�.���an�v�����k:J�nظw�D� �d�R��b^K�Ɉ=�@�HJ=%���hK!���T��'���9�I�\�o���3X�ѿ���t��A����D7,d��7�ڿ�/oG�3������t�������DST�`�G�����,˶ӳXa����*�^h�����n��,�rG��K�^�ʤI�"}m)� ~YL�N�b�Iҿ�l��p��OgX :`�I��Z�kSѱ���N{	���)L"�U1N�����Q�������Q4�d�� ��B�s�Rq��x���R�20y�Btx��m*{0F�Rڅ5��Sm�4u�j"��j�e�OЧ�\��,[���0m"��̀�^7%�*�!�i��7_�lO�{�!�¬ ���rШ�<by�2QH#�,�5����ߕQ�/��+��m�8L�� �����?�[#�'�u�����~��0TN�loS����$��&N��ԁy����#��M���}01� ���̏,����h��(tV 9;�pdׂ��%��Md��pR~8��[���&:��jP�Z���lμ�b�x&H���`|pU�)#_�!��Սm2N?u�\��K]W�c�˂dg�Ɩ���V���]���'ؤ p���~��5]e;O��	�!A�s-Y�P��%\��V>��ޘW�'{g�(�w,�L$�Nة�}�駇}�&�Ű�\g먑�;>�O�E#��g��1��x�����l�U�k��I���5���0��̋􎷰�V[i��Azh�1�Ig0���Т�#T?���#���C2��|Ȭ4
�2[ak٣��~*�����a��t/}9�?��Q��.iZ��=�� �c6�ղd�Z<�ֵm�l	����&��b�L��?�} oQ��A��^>�U�9,%Z�5��5�F����j�� �Ct7��^��Q�5�n��a�^B�RfM�±"���Uq�_�+��	;�Q�Fs�XZr����/� _�B>
c������n~!�N�t�]G����}�y�S�7��ͅ!��W�<�L|4��`>,l�S��پ����u��{nb1{�t�p��8� J��d&"~/��F����$k��.����tZ��O��	Ql9�SX�q��mR(�q.���K��)-far~�i�IKM�U�NM�(QA�b 7p�]���M�.���H�o��}��K��}�Tj%��{�� �@3^���{bvx�T�I�Xz�-ܣȀK�(
K�PZ%�(�F�異&}���̅�x��)��q)&"0�pO�h#�"�1FI�-_0�,=�,�)��'��QFm4.�*h�H��2$�q���.h�>0Q�(��$h/vc3�W�E�TR�Jب�_�Α��`Jx�*��=�8��;�
�����������_[����L"z��_��>D*�#ك~�C�f�ypd?�r>pA~��mgZ蟴�6�L1��tp�R�fA֥`�FqN)9,��Z��-�:��z$�/u������;TB��`�L���t�\�e;q~� `�/4�X�
��Կr6�(����*� �:�%Cr����ӛ-D3��!�g�4���5?͍�c@�f�㵐?�j�:/�k��ֹ�W��<�(�y�E�n�����������)S��j~��t��+�!�
��:�)g�k�� ������S����!�'�w&@rnUZe7�q0O�,��,)�+�;�t��\M.!��Q���7�a�>Y%p��@3��p��v`?ҷ��h*�w��SWj��˟P����cyv�%���q"�÷���N�t����@E�mZ�I�0	��vso<��!�m� iE>� t. �nݚe�u�X����|)��g�B���;���m������b=Nޅ�{�F����A����Ѩ\k5�8�#X�g�ɇ>y��Tz-m���ɾ2� qG�u|�gc�
��:Hç��a.��*�-�v1e /ۧV�ghTw�6��D	��ѻ���JV���<�V�I���<Q}������#�z�C1��?��{����'�b�Ǭ[1�\T!V�j0�vg�:F1o�&�@|���v-�&��G��Xa�;,��[��':��w��)� AphbFMS��D�+���m�͇3F!�M�R-��*J!~P��P.-F�w	�!>tNg5X����!dT��=�5 ���=��Y�~{��;�)���SWn��]`!`%�����i�|�|<��=��+BX{D���?
fn����
�1U�lly+�Q^A��@�ˀ{��1�`�#X���Y�K���Y�x����h� CS�6�p�r<��q�8X�WI��z�s�QH�C���H<����ݥͶ�0c�%��<��m;	#�Bg�gZ%K'j)1��F�:-W��=�& ����{�؊��^k�s7v�V_.ݗ1k2�g"���&нOú\�� Z,��7��
��YJث	�T�����8�\��m���{�s��5e��QD�-`v -i��[t��Щ���sO( ���|�f�|?�N^a;��� r-��Đh1"#uУx�V&�t�y�������3���ɜD���u4a.��\m *��:�N�}b�B�T��?�R܄�n?��͋����Ѧl:�2��{����Ѕ�=�M�Y�� ���F��T
3�k=�!�R�Q�}�f���d�Y�m�@~M�WM`'N��A�n>�&R7��!��S��j8n�Z��ٌ�����s��n� 8ᾮ��5-w���h����XI��Oq5��n�*��p7-ż9t�9X��Q0�1��$��Ǳ]/�;����j�n� y3d,�~c_����F#������NDYsWz������|����iVr|�G��^^1�g��w!���]�_v0l1W���-���8-LQ�E�U�������3�Ύ΢T#�PJ@\-;���x�7,���S:��.3�	����X�{��$ ��*r����|4�������;���O����C&<a�~5����!�/	RR���S0��5��:@W�4r����T���� �EyWCSC)��v��l)�L:�A�;M��y=mct��Y�3��&�m�p��S���bm��M�ǔw̞�}ʤ�~l��@�����֢K&q��f�ŃX-�L�֠�Y�4�� ����MFj�rGy	TC@	�)v��TH��<�@}�{�@�$.�/IX,ܨo��-�)��Ҷ\�CJG>�O+9]�Ԓ��u0�_C�7W���dȴ���D�8�B�*4