��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U&�0P��Ҟ��G^ф[�+��Bq�II�� ���&D�7'�@�~�F��=�5��7�׬;jdJ�W^Zy+�ج��w1�N	�o/�ǽ�ab��/�N[D<$<u&<��AZXt��5|���w'�u���ʿqH%�z"S����=�n �K�@XC��'��N�����g������]��"�nc���&h`$\������z)�R�-�����`��,.�Q���5y�ng̽�'�r������Ƒ�vMP���*�(��c�L|���������V92t�:�L�7`�سZ{���9o�F	%Dբ��I�Q@�Ć��(R_�}�jBD1rx2� ��Ct�ꃮԲ�!����0�sY���.���J�2�F�,j�Z�6�p2p^F�@�;>ѹ#W�\s��}r���ղ+��{�Gt\G��w�Oꤠ7
L�fۗ*��*����D���Z�q�M!�!@5]���L?�}��L��0q��Im�>���'
K�pRϲ����������0oQ�;˩���
->r�+$m��	���5.P�GOO6��"��
��Qᒶ�9V芁x
i)5b��<����Y�C$"�]���(��yD)�z�D�ߌehwp.�����)��l�s�.pZ�Q~�m>��_Fj�{�E���j;hI�����zB���V�71?��_�,J������k�R};*��V��i�[��	�<Ԫ�x�ƳMH�l֕.���A�<_^����OX�~`Rvv�.��
*b���i,�K_�}?:͍��g�����N	I�
z����ڻ�����f��۫���Y�o�H5��x�썂�2��BS�Wx��B�!�����q�`�T�����M�8i�o6�oƱ�����-mm��|��ҕ�[�j}����4d|��B�ox�v���U��	��,!�K���~g�H�@G��:U&w�Ø��� &�'�J��[rl��K>qC�
_H�I�Υ�2��|�����ӧ(�w�H����:%�E�¦!�w8p��^R�k�ڟ��V��|L�k��X�	�Ԫ�4U����=�+N�S�H�v�Oxb���d.��Ic���8�mgs�3U���x�����&�h�5h�c����|�����|s��E��7��VN�l�h�V�Ы��cB淦"�`�XY<�g��~���;���`��)`g<�h��È�)L"!ܳ��T�̬F���o�S��'�?�ی|\Ċ�nf�RD��[��Q�%_�-24�I���R�ȅC1T��*
��AIr����yJV+꟬SV]�bQ��:|��Iٝv-�����Y���$a���,�.V���S{�'!��
L�1U�Pu>�G����d�K�Qg�o��޼ۀw�^`�t��㿵=�����y�;�K��H@%���������^@l�֜r4"�:�$��L��_��[WC��C��p���\&�Bȋ*�����Y�����L��14�
�8�-����D�pP�p4��olj����{q|���O��*�Ճ�.���t d�z��FR�11W$$|ň��.� �g�[����7�4bY�+O�
1i�`�|%fkIe�Z��b���w�-�W�}ђ�����í�-}����7�M,S���}3N�Vδ>��=*$��s��Eew�
�_�}p���na�9�	Hj��m��[k%��?�T�{�ym���$�g�'��3"D�]D��?Zn2�����ϑ"R��s����������Ri��u{{�0��8�'�h��ڒ.6�帞�1�~p�h���+���m�"�*��t:s�����M���P!;p(��Ǫ�B/��oE�JK%p���	UOf9N���4���/��,��ݿh����[3=XF����DpLu(��%�2�uS�s�����	�,:��G��j���3�5���K �c&��9�ԉ�xwQ�>�jLOVc't�R�,;�$����)Jzuo�U����)���6�o$K�������	��l�#��#��!�W�DD;ᵴ6T*����Y��
8�r��ݢ�4���/(��?�	�C�d�+ T��u��pF����E�L�Mؓ%�\�l�>L��%Iצ�#�N����F�{hqr݇.Ғ�PVJ�H��jI��'A��X��,�ߘ2V`��-��a�=���C(ܹ���QqMli�~�����ܯ�������@^�Q�i.%60�������>�c7�W�����0Ex�}�e #���E:<䪎Qe�r���FY�J����x�ǅt����-���O��}�Mi�P)����"��ߝh�����g:���M���Ȧ&Z{�m����j+�t"��x�'N�~BI�{}�#��[_�:��32=�b,��MBo�(�i�
(F	�"TFX$�q����
5�t\r���j�u�NlÊ)�LX��������_�I1�V51��O���K�V{8�M�Oے�C�˰�_���L��hQA�m��Õ^a+�oꋛs�}�=I	?f����ݽ��6T�I�KF;����0��K`���
%\��[͜�(�g��isY�n����[}����>è�_
�#��HBtTJ��)+�v�ڌ���i{b K�v��s�ˆ����GɚmS�;�2��8�E�䯀�� � >��i�,q+Ӿ~�vj��f���O��8�K�q�ǃ���Ob���S��/o��H �)m-_�ǋ�����"Z[��Ea�8c��d�Z5�z�	��ڻ����L�
9�hx���DT��6����ō�-����C<]3!�Ù)S
�zP�n��J��߂�c_h���c�nU�F0i��4W�.c�;�� ��Z>n5�/�$��L���2)e���|���Ȣgأ*eěO '���ƽ�B���Y����tB�uLݤ�� �Z<���N!`fW�k�a��5BMI򓓚�b�8[��B���F��H��UzM�<�*�u�y�L�5Ո�X��ޫ�AEAJ���������B$n;e�2�T�s�"ܳ"2��`�������of4�'�s|�cwv�˻ǅ�|�k�cNe�j�P,W��h_>�j
�]� ��O��<-�#���)vuev�-��(x�4����s�X��Z��@1?���Fx_Ct��y%�k�y⽿^6�%�^�wnR馨�X0lV�ǿ$Ӏ�y9e�L��j���w�4��2�🍈��H����'�O�|Z�ՅV��<��6�\I��4�i�O\��p{T���s\A�d�JΆ��H l|�:
��TP�A� ��(j�*�	���v�X"�T�~�������}�\N���n�|�KpHE��S�]H�CW!	��Y��P}����V%�$�5s@�b���X�<�XAh�\#�#ƭB�8����A6�.�Ip�:��9�ɕ�}ہez�� V_?c7���eH3͓�3,f";���9�G�������+{��*����l�7y�ET�
�p3������T)�y�W�`h��uV.�y�ƓA�/	���M��G��p%�&��&_B-[e�o���?fj�_�^VL!Y(�<���� �S���(NF�N�iؒ��W1n�)!�h�`��rJ�J0�?�;��4�(|g���Uڐ���4�ɱ��q���x4���L��dNY�