��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5��·t����O�ihY�p�[��s��o�C�>1�M}]s��UN�[6�0>��r�W�Z�5e�݀�Ew,b!Ə��8h�Q�ž��0_�=��('nE���i܅Ǌ�l�T'�j�z:���ѡz?��@?�hZV��X��D\���52�ޤ���5l/PEp)*��K8������W��䗰���.
`Ed�+֐�L��E֫L��Lw1��W�b�8%,��V*gH�tB))��Ԛ����k]���,4H^�EM���/vܵ~y��ӶZ�I	�p����`3 �=~XFI��=���)�ShfK���aA]i�?�IG��9�a�Q�5�.�z-��i��k��7xc�7�hǼ>�!r/����e��'S\B8ا�긕iI�5����5WW�6,� j��:7(L�	��?#���%iG��q��Δyox���?^��A���c�>����9��g�ZĄ�3��ʱQ3�HHEҶM��g,wq�GmSpoT����D.`��i�lT�Z�#� #{�=?AL󮡽˧n��g�v�B��s��*L3�����Νwp�+L�(R���[l^~���`e����߱�z��� ��>#8jZP橿,��]� �(���2T�\oG^��o!�_�ۏ��Q��ѲXp�����:Qh�0��̋KA�D�g/�OUO[�\I'����st���1l��1L�6?�l�0��3D���ǐE�(�5_N%s		;1�3��6cf�p������ό<p�H���V>�3F��^�7*�kEDEV���~[�q��!�*�i[_�H��_��a�p�\���l ����,�Sh15�i�!
+�i�=E��&(`s���S�sz�B�(�k�GԖ�C,U�1����O�?qD��o�:Iǭ:e�'�r�8��CO��b�B�^��Rh�h~��b\GT�'���6��]x���S��Z?�K
�ݬj�HM&���x�xX�ځ�" bK��"���ȃ�:N�R#AB�ub�!|�9����C��HZK*����j���FQ'Sa�'��1���YM�\}�N��ţ�6QSQ���	&���l�}�e��p���)BI��m��*�,DzR
W�D��K����r�#�P9��0囔�O�w/����)�M�^pA"� �{n�C��û>���:�/��bbg
lz�	�?(�X���w�F0+�Y�s�Q�~V	�kjAb��:F��P|N�d!�r�,�haƞ�3�3�Fd�Y�V��!}��re�&XvP��*���N1�ε`��6�%y� ��k<�ʒ�jR*����`|G�2\{�L;+�o��p&�q��v�-$�"�Y�T��6����$�8�:���0(t}�!
�Z`a�ئ�bKce^�n�L�tr�);G��-L�c�'�f�X	&�q#'�$����(jkb�H�WD��^�7Y��N2��E.s
���S9�J6����F��j�.bX�g�2�\���a"u��쎺F2��M��kMO�����L鮥��\���u��ͨ@{2ke�D18��up�r�Ӆ��k���ZK�LV|f�P�*��*�����.�[�W�}�kѧ���Pp�^�����Z>�p0�.��yu�J���;ɿt^Tܐ�ЈH�+1V�(;�����x�������^�u݀3�4Ò�T�0���ju�7�HN���»��a�������]��N�z�󁓘t#��#~N;]~���d���P+6h��2?���/���uﱨsb&*F�b�"��?� �: ��iP}��=u)Ի�2�GsL1l�r��bE�P\����I�d��IYXi��4ٵ���Ύ�������oN*���m�N Or�8]}�F�<�I�������ɎR�� ��9i�1z̧��jF@X��H8��tn ��e�H��/oچg7��Q�ՅhQ��� �]5������W��ޔ����V&~G���(L�pX�Fz
���ލ��X%6������L����(.��%l�[+�p�;�����8D7G�qV��� r�rP�c	���zs�1�eg7��U!��eǤ2�=�h:�R�BH4�~,� ��,�q�7�p�T�Eoy�R�ߖt(�+�]'��Ai�6�	5��\�4�l��u܌*:�S�޵�n�nrcR�D ����V��~n� s�*��.uuJ�D�?̮\}�h�:D� �(J�����(-����&��ޥ���Z��~�v�˅z��(ύ�ljy� �p�R+*�A�	��Jz|�'�Wt��Ǚ���5�&cO>Y�8�<N7�L�����^��}
��&�E�����&j���$_��kCpl���F̜5��(jv�.��JJ�g����\�4j���I�NT�콜(%�}k�)� Q5��Ej��Nu*>JZX��nS�6H�JK�����p�S��Ss��@���cj>٢�����y�u�V� 6�5/�����!����Zj�+/))����
gFx�3��֏g�~gϨ-��jn=A��B)�K�8��T���ӣ9���_~��)[c�ձ���U�%��ڵ���X}p#�X��%i�
�r����i��I�_����E�<�3�G p�Y��r54�M�[���d�!���%�-{R��M����@3�S/��� �;���7��k54��qv��ŌA�P͠��c��a. u4h���t�