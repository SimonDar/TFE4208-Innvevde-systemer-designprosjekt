��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~�f�?|�ў.mh� M_)�U���l�8��:̜uYs�O�ƫ��<^Ƅ*�Æ+D���/�̳�^g�!�U���`���ע��K�`���gҬ��M!��fp┿�;a�s���{����T6��e��B��jG��r+�kdk�I�[��1��<O������4J8HZ�Á���}�8.�*`I{��EP�H�����L���T%x��/���Q��n��1Z&�v�W��I�7QӞ���e1�
w�1A"�l�3'�4%�!���zNU@j�'��$��/c�G�I$Ν~q�P��'���>m�P�2<L��qov��q/`X�����?w`���15e��-H��Nr���Hsk�3F�E�l��8>�+Ip1]�q�5���H ��c�1t�R9�k�)�{�`*k������3tlz�@��wm�$�IP,���Z�~;��XY6����^��ly���3�ٟ)!Vض���9���C	����0܄�8�o���!ӄ��7e�|�la�]@��cB, ��TdP��EϾUj�u	'�#ࣾǱÜ��uKFG�?����8�����Tv�.�{f���d[��R�"~޺��:��3yM��gFF˯�Ա��'+��E��~pծKe̛&����DIÌ��L����2�~7qN�$Eg��	���?�U��)�2)�~8��ݰ�
o����3��y^��Nx�FK��E�v�l��KM���T��Y30����>��Ii<�� � ���*�d��4s@2���$�7z`O�L��*Pd����^�yF[���1���;&;��G�&�R�V�|dܾ��'�>D��X$}��wN�6Q}lq�}C�09q���$t����~��P��u�Y��<,��礥�����ς�*U�w�~T6�6!�Rl��\�g�1��GS���;y"�/��������坦��[�؍-��qr�����?l����͛��dϺF��:a�G9�r)S!Jy̗�Y�/�Wv�B�1:Q����15#;+���/Ì�Lt*#��Hxڂk�g�{ݘ��L=�z�n�k螣H��)�Q��pu�i�N+C��"���ߙ :��C��Ѫ�>q����қP��gڰ�?36�|��}�ph�
~�%�G0�;T(��ٓT�QPC���>�@�����,��-\d�;��Zv����јq��r��;���m[n��l4}f����7���E��ĽbS�����ZA+����6��+�uB���`xh��j%~a��C��L˙��O8�*�RJA-şi�/�m��]]�&�B����V���v�5Q��5�62�V 4s�����\���Y`�VN����dL��P�#;�f�����K7~��_�ru��:�z�u���`�Rԏ	�M��Q�}��<Y��{��`f��FU�,������Vd:����t,/ ^݆�<���e{z@2}�l�M�������7v��~�b�1�^ᦑ)���];�"���}��0�($;j,BS�il��X!�'ɽ
�wz��u����mh�}e�� :D3F%��_��/c|/��\�TM^��I��ܣ";�ZK�$!o�Q�����Er6������s�aPm��n.�Wl%(�%���tؙ��P��H#tA� #0U츞D'��a�_����.��������ɡW��?2l�	QHsF��c�ll��m�P�)k���%`s%\Cאsx-�2R�?��(
�>.-�ҍ��,|t���C������4��_��)l�f�2ѝ=����!�v�ȼ{f�K8�mkK%26K��5g�TbW�'��e��+y 0R +{�L���+�R�R���ڠ�)��q���m�_|F:E��0�y��q9�[m%D�o*:�d��A��!"p����@}��X�9�'���#�.
�G�<O{�����c#���x�/�a���ަ��k���8r�~���"���Nw��J��9����赃6K�_?[�ѲH��&Ql��߀�v�[�g�&���2��),�������kP�o�����f����+���~!�նBo	��u�ֆ�"�f��iW~\�)f{`�o=*�3#�^�n!Q�`��6oDg޼���sR��1�%�6���9���H���^c1�~��7=����X��E:-��ÿT��2q���i��%����6"��/��<R|mvTL��ȳ*�g��rOhg��v$��{R��h�iz�e��r�Y�g^�:R����-U�j�c�X�<�{yu=o�Z\gDgS0`Q'#P�Y:Sb�؊��\��������2�3)\�\tb���}��rJlw������å�2���ƨ1��Y�}��9����L{���0d�K��{�4�h�9�\�"8|�2�S�3ͪ$����]�f��h���������&���Y8⮷ߛ(-8���~ ղ8��.�#>cA>�S��7�*��4�>���k��Jq�Z�Xɮ��K� mX �{ռH�ǸB|�QC)9OvM2�ؓ�AB�D���#`q��"�a�2�l�B���5�Z��A��L�J��c�)J~c��X_<y�lt́<�r�ju���]���S��R;
�ѻOmAa8�E�V���.���$Ղџ*?1ZƘ&��e]' �OQ��u���̃;�C��F��I0���0!t��>�D� ���y �3�`D��a��'%��V����z�������΍`�ů�B"
5A_H�{�Jhd5�����Hr� �̿ ��דZ&��.���:��a��Y7�E۔AxQ�"_��J�j"PWf�G��qA�T��䄻�{���-��������s�ﾃEԍߤի��t�TW�Fr���|�0����~�R��F��v�Bjw�Uwxy�����=�%F�{V0iK����V%}o2���l_-�w@.
��uh��C;� m��)Ķ�#������W��?��/ⴑV�J�q~D�W,��
����y�����h�;S̓Φ={^�y������0-� �B����!&b8wl2�W�O�*6^��1nQ�Q���q��$� Q����C����و� �ΰ�2�9���0��&���$E?j62BQ�X��C
)�!�uh�����������yT�x���)e��m�Y���;L�W���]TWA]U�Y}Ԟ	S�����H.�����ܬ�H�C������B�0��_Cg]�8M��+��2YBQ��|0�/��r�<�"���_\v�cS�΀�h;q>WM�)
y5�O�����>��N������S�>�H�K ��-��>½J�}��½.5z¿4��wPu~X8M�ً�1|L���QШ����{�͗��{Vę�l��;c����2Q���e;�*����y��)�$�{��[b\�!xDO���|pWd��ň�����~�!��ӏ�J�ۓ,h��(���y6��M�PeyfG�8\�����[,�����k��H�ڮ^��qSQ�Ȭ�f�xH���Ad=����i+����ʕ���nr&���P���0ZS�[���+Lq�>�כ��K�oUx)'�P[~.�=�OʋL�]��q[�h���B��O2���.,�z��R�d��-�F����{��7g��F�!�Fؘ!��������Z<�-��<$����)�e�n9�ٮB���C�Wŗ�Ρ�yۏ�j��A��Ĕx�e�&3ٓ�L���Z.�3w�Am$�>b��8(]"z��&��6�EϷ�����N�N�
J��NuほMe�Ow%����ڣ͋r���ێ��������u�1���t�>n8j�]O�@��63"��9->��?��(��\b�ɱT�D`���+�XJ��*J$�@Pww��A��1�f�N���;���k=��P��܌��V���k�$lK��,ݪ&7<2Ѝt�.�0Tq)Lv.>���L��<D���J���9�'fɣ�,����������'�Y[������h�]��{�G)��Z��6M��~�q���8(�r�Lݕ/�Hk�"\�J1s�4�C��(�M}��;~��X�d���rB�3͡"���ԯ�Xrn�'�=3ĳ#����gX۾�g9?�5(��+4d�~1���!mX�Ђ֏	J9}ק2̏Hm�w���y��{�����T\@���%�~1)�*N�pG��N�T�Sg�8��8�t� ��贛��~0k�
� ϐ���V���ʜЃ�$b6�P8B����i�nͳ�&=�)j"]��̯����p� x;��5L�o_�{�j`��M2c{�-����x��5ި^fa��$w�'$ض��]�]g����<��l�6�ĥ
����JG`�ǳ!w�DL�f��)S�x�o���B��-�����}}�?�x��͎��������,��}L)1b5-�Ob�/i�Y�`ӛ@�Q4����0���نr6��Fim��^f�r؆�~�H��;}�����i�N�RJ�\��=�� H������l����+���L(�+C��g����tv����`��Fp"�?B$�h	�����!:w�#D��l�KY�.X�@v�-�~��}o�j����K�;�k=v5�"{I�a�k�g) �
�֕a�J;8UR�p���6��u#i��Yf���#�fH�:�N���8��_Ey�ﵧ1�9�.'x�pҍ�
sn��*��;������RӺ̽��@�@^-�s�!�w!��c=w9aѓ(�q�f�*V0-)H8&V���<�r������9D�3G�:-N�8�e|��ĝɅf�2�����⎚�n�W�*�� �b�n
��SGq0k\o|�mS��彑m�T�����w�SŖ���|
�]����$ 
�E��I�zL.!0ͺ:�����@y�ɞ��_9����pl���?j��C/w �Q��;���!��M@d-�G�od�o������#��ou����^��!@X��5H9�za?ΎJ��o%��$����d�$z�%ۧ���	��C��at�K�?;�G�{��tP��	��v���bk�P?M��\W�q�t<K-�{�o�����+���q(?��
���j��݀$CD{y��ԉB^SzBGQ��)���fZ��U����Tn�j������Z��En�C>��N��Iu��7�{�(���K�����%�+G�e_<v�'�g��DO�{��V���ON�D�`P�����$a|Xԙ=�W�̉V���j�j?6��I麯F^';���w�Z������M���\�z�W}�7�<����2-����	��ɳm����m2��	�y��b���e�ۆu��[��o1�� ��u�H�J�V#����
3��^��M���q����H���5Q�ȭ�R�DOw�T��\���<�@����ё�3Y�nؾ�r.��ܐ14Z��TI�Ef�L����Ҳ�w����D,s��_�#Q��<en�����XD�0�B�R4�v(y1	�K��9��GW�l$�@�c+~n��"�,�Ҧ�Tp�5������i@ބS+󿗬�Gw�wO� �԰����@d���kT���7��qD?!vz]E��`��E�!<�b��S ��%��sʼ^�.�j��7Q��rw$_��4}��N��apՀ�E�
�)�e�7|�@��k��'n�� HIq�b�?JIK>�p"�{�YC����GoyJ*�GK����*J�  �ZO�ǟj�TЅ�Z��o�H��2�Ռ��r��g��k�Z�uz7�n�R������ =��cnM���8�oX�ye.@���ۖ�D���[�N$�S�me�F4L�I !�9&5�(8���i�����&i\h~O样Վ�yzɫ���
 �ap$����{���P7$2��*�H1<C;a`tmMN�v��#ǃ��V|@Q/i�<�6wo�?��&��/-*o�m�V,�N�5%��1�w��&<��y��zN�/��O�w�I%T�-�AoVc�:x)�~��!so�E7�oq>��'�y��\��i����I�p�@�[!K����B�K�t'Is�\�*��4ޮ�p}���	�}Q�q�������5��l^,��S��ȯ��s�F͠h
`b��V���p����lZ�l�� 8���u����y�����s���o�؟��O�%n�oh�Na�f�d4)���f�W\�����Xj5�K��1c�Y3�̓�8�Y���p�n1����&W�����W���]7��,��(��t��H��Б�h��Y�S�� �:yOS�]�`Բcs��6u�����YN~��Bv�pzs$�G�魲�ٳ�>�tj�XLR�O�����P�F7�>cܽP�;f.�BNI��-�6[ɇ������Ef�]ɞ�k�p�Y�kg[zk(v��Lb���de�&�$s�S��Dʽj@��9X�.��U�{�j��v)`�#Y�n27e������?��չr��W��UB�v�ʂV9<~��줡�~�q�k�}6̗���5TQC��=����T���n�����s������ݷifaE��%Uh˽��&�]Q��<���1�>k����"O��C��ٹ�#��os��z�4Ě�<�-�:~0ʳöۤq��Z�fV��0��)(��v~�����w)U���e�b�L	����Va�ߩ�����/��K�??&L|�'Un�&�9�>�αLi��KT����LB��TC~X�?����EU013͚N>�35�L�Kρ�d�����У
B��O�؁x�D��*n��)�]�//Z��nK&ALL'{�.�3����}�B�s[��7G�l�ߎ����_��h,P'��>=Z)SD'��{?F����M5���c��Tܧ�08+�`���5FOZ�cWw7�W#�fr	QI֢���G���6:��/|ș��]7�d�w9�b�aT�G���:�4V�g��qD����4�бɫe�}�kؕs�t� v2��	h~ሎ�{��(#ь��ƹ��QE���L�lΐI�q�G/Ai�U<���2LSu	�:�wM�F�,y��(X	�硧:�g�l��˖��`8�	�9���i�,@_��t�2��hsR�w����w�������=���w˯Ů��#���*�@hΒ��ۀ���������V�p��ढv�Ra�87?P��x�)�V~!�Q3�j5�ޥv��_V��M�|M��s�	�C�Kr���u.C1C���2gJ�]���eU�;������p/A%U�Jj��I��A�����^)gD��Me.�����t.*fK�T8�oGm� SL'���o��5l���_�#ɧk>p�Y"�N!ɥ�͚y������(a��ˢ!�A�j�4hק���*"bycC+�G�"%�����27�Sz"��,��-%�|eX�fD�x̩�/�b�m���Qϡ�-����HX����G�DC�VxzG��R�b�H�bS�IKQ5D[����<YA�{f��&d�V�U�%�f�T5p�(�+�U��n1�=+3�E�qr�"ox���SQ=�"S�3C��XԅU�/�]�|"�0�a�d¹OvB�/=,��eł��D�`�eF��,���2�.-|�$�D%갔��Iܫ�Ma���;�����x� =����&Y��ܰ@�n� '�6F�K�- ��>oH!O$-���P���'G��Mz$s�h���d����?��Z�U�E��1���9E�vZ���$A���P��Wߓ���	���.> 03WC,��W�����^�2.�d���%ݡ/�4�*e��0	�6,�r���0p����g��&�l&y�|�k��io�Pi+U���]kLWn�m75:X�W��c���rh���8���/ք�?��m�3�2�;�����7R�މ��K*{���㐔���8�Z�;tB& C�I�6�'���J6v���LreQ�`��1���g��L`�\��E�*⁘�uR�o|�����QK��R���������,l1�UC�)�p�Hl��G�Hg�30����l/-i{F���;����E-�}Y�6ұ	i!����O�Rw%J���IO�|���{�tI|��&e)r�5���;��C�� OΊ_�ք����! a�
L�U 
>���MZ	P͸��n�L��Wu�����j���B�Z�2G:3�g5<��Ep�y�آ#�����@�Q���o{_t���P�H��Ř�\�o���&���1%�.�?7P���e&�@R��'}�y?��^}� :�$���T����:���|pȇ��z�N�[9� �*�q]ºr�hP� �t?CVZW/���,�%�mFS�t���2���S>WJ��]��ieY¬�W.?��{���E�N�$���8�O�Mv��^�n�-�����֛�IYE���LG�jh �h�xaD-�� �aN"�ܞ_Pf���N�4�#����<��r~�~�	��	
��J�8���/j�wxx� q76�uꉴ�u����p��ΊB2�s4����+��5/�W��ɀ6�퐄;��qG�����?�&v�-ۛd��$s�YK��fj#�FD�
Sq�Rv�~��71����r��G��>g�D������֭�n^H��`fD��D���O��C�6�F�ӬD�	I}�E%\�:}�?C�=����nN㢺�� 9�鋘JBɝ��� ��@��6aޚ�{S�1w}��	�OKz��"����+[�|�v�*$���脴KI\-6B,8z�G-�aЊ��O4&���C��3�I&ba��4�T��p:��˨z��5��P����e.#�<e�퓢g5�B&�+2(�R?K
�6�L}7��}�ߧ$v-�"C, C*�Q�+��"��$��}�m���{��Tb�4E]�Lǫ<�ܹ��j��2�;퇻Ի�����c������_����*��d��h\��h���V��J�G���|bƫih�L#���E����.��[2���ϕ6[L��\o�9t�HbI�9���rdA���('j�c���u�/��Q�p�y��F�8
�=ɰtGs�����t;a˩1/����ay����/(�� �eו���=�U�2D����L�/�$�����H��2;�
ù���7[j�~n���/�@��~�WO\���y��&6�-�\�95�L
��i']!_��}�z.)�W ~�I�:m�q���ID��$nkI�Md��9U
ļj,���8�{_^�����e�k�!��M_��7;��[Z�0;P����b؁w#V.e۞�8�4;�A�B�o_�݊?��� ���`�����)As�1Gg5��UB�Ņ��$��6{gA��D��9�㒛�!C�?��9v4Z��/�7tυl�Q����VDj ��f�Z� �:���E6�l!�2�0�'Sؼ���f�xU!�0r/��f���Z�@���(�$n�v+sR���������P���?w�_�㞐c�|B��x!��춵���+��sBuϬ�S]��k�֡}.Ga(�b�[��ڽ�<G{�ڄ�H,If�f�.]�8� �+��N�gU�O�I�Fb�D��T�����/��6 ��,_f(��;Ĝ7�1���:�����-˻Kz�ЉJl��jɤR�s�)�j��|����+�7>���k4@�,\hÿ���̸t�pA{1YA�*y�G��%����R�(���y�H�
�j��r�s?��\��E��QA2��.�heuA���Mܞ"�c1=�uM��G6V$��M^ğ���[i֥��`Y��3d�!v)P�g��wg��җ��+چ��]"hN)��ܜ�p]���b�4�>{?���f�0��督d�(���=��o�æ閨��ꮴ����qD�+��=�O���=I��W�z�b��s�]���K�$�EUt�|�`�5� �}���-�C�_ڛ|�w�A��fw��ľ��U�m��a�oc��R��E+���{�v�F1�M�.�_�y�7/9G�ż܀��{�O��c���������I�!p� �����������4�����2�rª�7S��Hv:%��ei�_[��#�[8X&�D�ps�!���qy�^t/Q�	�`�U�(���)��%�-ڂVop�7bʱ�!V��s��|�P�:u��)�<b�����5Z凉G����/�A�ӱ�����K��Ƥ���7Ν��G�������w�v��~=�����:�#���^0�=��q;f���Kf����;�����ں� u��z�g�\���`p��@�~���!���z�*�P󤑁=B	|��M���#�b��r�-�H?O�/e�h��3�")#_�܆���k��e˘Cg�ƿa��c#~����X���le7t� J ���2�\g8$�K.�F�|n�ݳ��D?����nM��a:;�5^Q�{q���7��"ņ���@�@��m����b�_���@�MQCr�q�8̽?�+���T��/�P '��k��̣�#���Cz�/pC~�`�{�����k��XNm�������$�_�#����⬷gLC)��y�5H��	�J���+�pS�$��+�
�<{��YN2�n�>B������ES	��>e�܉�w�	�/��><Ul�]��X���*��u�����M	(W#zߓ�Q���K�3��M{�3ǔr�G�\��/�Z}�PA��y�K`-N�E�-��߱hŎ�	X8��BpGc�8��>i\����)�<�".l>���gc���D>1IoiGA]��2֙*:�*����p<F,����6�b�YE.�����"���X�k�^���`�G�MC�M�n��vS���G}�� ���n�̡d;�tX�ASD?`��0k^-���q1{����O1p������B�������q�bN��*_��N�<v˫���X��)�8����*؞�j��5�A���3�sGP�OV8VH����>2\�q_�榼���
��tdȬJ�^"���5�cO&��GR�^w2���v�c[�Z)�8����8�9��@RZ�"��������l�1^��+x`L��a<�j��LE����82̙zߞ�`s�3G5�qS��J��E���",��͹Ie����#�R�UY$9��|�k6A�_�9 [�P�WxQ��:��`�E�U�D��������Ӊ<F�Kw����bX�Ї.�W�f|?�#{;��e.ɖ��
<�x[�ӱ6�fBR�;-;�!h�[�I��L�E*�y+	T��/������ӵ��H��`.]��R ��xLM�qW����nć�_w����S��B,ݸ�C.��Y�f�@�i�#f�*�%8��vW�Z��ޞ�t��xC<�v2,�b�O�j(����im���x�s|GL��lh~��
������==���}[���K~z��ݼB�Y����FI�Ѵ��\�$�)Z���Z���a�Hn�k��$9&�^=goN�R�ېj_@;�O���L{�9�7�ty�0�f��&r�<��c~���fj��H%#3��7�_���z�ؑ"��F��/�=��t6�wC��{oFy0��@�byJ������"̆�$�s���%q!���ܲ`���uA�1/�ՠU��O2��v�O��F�/�y�or~<9�o��
l�׼��Ks��<����z���V�P�e���}�U�t���d�hE�>Rpa�cU�ו�����r�c�C��V:�ƭ%��G1��\����ܹ��A�+��x���ݛ�"��O�AlDNdY/I�`#��t7*�~��(�?Ry:a݀�xAq����+�g�F��\�k�Y��n@�(~�����?�r$J�v�#��ڮsjC6r֛���G,��iٞ[����d��&d��~;pS�iդd��&*nɕ�o�rK|
��Tq܊��G�2����z��s���q+A�m#�ȅ��W�i�;x�Ɇ�1�x����lU龩l�d�T�󘴞Z@u�s;O��R<�iɚ(��<��<o1͍�&�SZ���*0�m_{�cέ���uC !./}l�LB��Az��`Ci�?���=��|�vf����H8hP~�.��d���=ƾ +ng�}��	,B�7�m;�FA6 ��=�)EHC���}nhi��J8�ܷ%�l6��vc�푃y㊿�O5{�D��͹���oN[�|f�˂��:�GF�ai"��`�V[L&A���>ZC������r:����G���h���]P]\���	����h�m!�O�}����3�g��s� GS��]��ӏ�B���-� y�b�YR��w&b�h2+>Xܳ��R��׮�^f�M�}�B��(mX�QF6@L%��n+oݗ2� �o`�y�"(W�,��,��G@��x4�kHL�[g��>�k�a�{�<_d��E)x��/�$%�$�i`��-�J�N��9?Ԉ���9F(�qxL�0�3u�<>���j���ކ!����+N�L�dL2w�� &��Q�b�z1����Z{��O�]R� �!��Ncc��Gy�|YO5nG.Q��;�q�r�8K�3��U<��%���#0����KTV���ѧ�z_�n]GN����$f��a��+�WQ��(�4�d��ڥ�S�����.�[�C0M�3^��з�c��}Nn��;(F>v�Z��*Kd:QZq-�̃�����-F1�f���.DaxI�SEx��ɭ2�n):w�O٨�Ud���dܒ:%��m�Xҡ��S��l?�o:�k�Ï�|}�`�u]�yK�k�\�D������g�2Z����P2/ݼ\R>Z3��>ɼ?MeOt�a'4��:�`��?呖
_����&�Í�=��;w��n
H�_�Vr�Tf>p.�v��/U�[yi">�̙���m%	a��R�-��1D�߽2#���/��-���>��x�g�{��aY����+�M��>9;8rn�? �jMV�-�c�,��<��8`�s_8ŵ�^��U�H�l�"�I�􈿮��qd��j� 
|e\���^�`[�����N(�eцQ�.�J��ؿ�lY�)&���!�72Y�ԅԯ�i��w�T;)I&4a���~�QQ�0ɐg��浝43��$�%�)�l�<⤵m�)�Ϻ\�;�e�u��HX����:f��ZΚJh|��'ߒ���'63��E �����@��J�FJ��i��ɱ�����5I���!5M��jW����7 ���etþj/��<B�IIR^!y�,��rS�4d:9��C>�d@f:W7�ɷ썹�5`o�v���H����+:�ߧ��y�?�K��g�;�e��'r����z(��r��e4$sf;5��2h�R�Qt"�*�ٱ|ܛj���G0���� ��ӡ�����Ը��}#��:��I�>�K���_u��d�������'3Рm5��L���/�N��g;��]������I��f��&�$�Q<g�mF<��/��ȚX7�2����y2���ȯ���06 �l�ˬp�ןCA޿�]̴��Zw�77k�.U��*�҄��T"1z,͈���U��s�%QZ���;~�kr����B��i�6LN=�5���6�������/�c
�� i)U����$&R{�4n�r�u���b���B���"$���ʂ��-Q[�G�M�g8�[�ۨ*C��:�X�}�!���eTl1�zmG���9��*���c�R)�/TfS�� ��uّ�,EwMI�%5���$9�cK��l�����u�^YDL��Y����@=����!,��]Ӗ���0z��WPu�XL�����b�^r2վ۔��JOkDd�/���l����Bȫ6�E�N8X9R����
���V�~y{�G�H��/?\Ś>"jM:^p��¯�i��LH!��v�L��Pf-�ш1��;�,�H<��k����"W�	���x�fe$z�^4���ak�|��4�g)FS����"� 
�%��K\�w�e���e�ňs�5��@�\��c���Ǡ��ך���΍�b��%9��BC�mNծ��0K!�9���Yn��{���&��=�mB�j�S�&���]�(��B���9r��2�����ʄ��=�_Xʱ���XC���&�/��>�U<!��m+�v���̖QU�^J׈<�Ђ�R�~���-�R���rW���ų��H���c�Bi��]05:����El�A[���X��0ެv�q��/���W�%K����L,ѮΊ���d��&d-�2��`�Me/5��	�� MN*�Sù![��h�,�
X��/cO�-���[T8ؓh�<(ߢۑ��J%�;�� �:�ܿ˯�ۥ������}W���ꗋi|��z}�۰�E�l�t�F���!�u�h�p�g`�*�Gv�:�A����NDD">�X'��6���d�l᫛� ����/<T4�K"�������
B�
A�I���ֲR@�������7�;���XN��Y�[~@�Cns�H�
	>�J��!��j
���G*���=eQ˝���Xt�ڎ�2��/ѝS]��p��<jW_9�@�d�Q��)�ը|y{��A%�fO6H�!�lT�e��)d=��?�Χ4�an�{����:͎,> ����C�̃�3"��t6:fD��$�g����`3v+^j�d%K��t�˒��Z	Z�&ɳ��R�MT
�/�5@�h��&���%��a�j�|*ۓ��Sχ�?ܙ9ËY��s��|ɷg�['�ԡ�E�v��郚#�xl	ś'���b�՗:f%'�&�����Q��YG ��|�砇\�����/���`;<�?E��R�;�|��l��Fv�E��Lh@P�J=�Iý�U$*q�Ir�1%�U\�6OPa���q�cC
H	�g�6 %^QM����E�������I�?����#�f���$k����u���ҧ���*���B���k9��v�s-��Z��!�P����'O��;/p	���о[V�����OL��L(��%J�Д��{r�j�78#S: >��� �G�* �^�ߌ�!�!l=�	����gU�Wא"�D�� t���R�K� �g�4wsP� ozR������7��4��G�-�\'=��9K����} ��*�5�nHF�U_FX����
g�;�0F�pM��Ֆ�q����e���� +:���D�zc��q��c��ʃ<շP�M�n�w�j�s��D��ޑz�_�ǷV�ts�W�¸��~��& GDDּ�C"������i��t����r�OiT	�B�� �vk���F�#����2���܉�]�a�f�>[Te2�T�C?�j�!�^Q��o���F��uo9��y!����@% q������p.s�+q�>�؍���<'���І]�]RcIp�e�g�쳔g�y��3������]Z��3a 0@�ΰ|�ŧ2��h.�);>���m��6�D�����T���!UCŌ�عY`��F#|��o�3��O}U%\�KC�0>��>�1&+0�?�z�\�m�z?rHB���O�[�.L�u�o)ֈh���{��KI0$�(p��ʸ�!r�:���	a�.���8�bVV