��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~	U�_K�-����(�谝�of00�,�#ʵ�r�d���(��Ҙ�C���FV\NF=�:ŭ��$A�b��q���@��@ZƦ*����VEĄ�F�3��cd�����Cw��Ҵ`��ok���а�a�����=�#7�M��� �� pa��w_��6 ɘ���a����$p�$���.�<^�MA��@�g(���:�WgSfWH佞j���z���V�A�N��1 ��к�5��
�B�+����m(YX~�Ƶ��M��v�_��suU)b���]��y� d����1��L ��v�g��JIB�C��vI��;J)��4��)��q|U�:�"z�j�L�����Y��3�
��Q��q~���[J�M����8<�l�ʰ��8���H:h�w7f`�Ƈ�Q5����Ѿ��T�F{��N�B/~��^�}<��[��N!Yh�!�UY8
��`mT�I�����x�s�7i�mx� 2�g?�z�6�[Ã�%�3�l�����f�/P傶0�D}4�Wm��������*u��J�⢈9�>9j���	��* h�T�Hi�m� �	�c[�?���Ok�bLX���_c�lO��s��	��������ac�uM33�Y���<�i��T.���T"�����z��Z�u6];��b"l��s�F�'�uu=��[�v�=ErE���'}sZ]��,�*dd�42���ĵ�#�;��(�����T`��W��/}�f-�S���F[�nx��`L}:��p[E��Z;#�fM�Ƙ��kMY����~ׂM~u?g��Y�=�.���<�L�7]83���^
�����Ň�}��2.-~b�tz���-�<���Ve3�o�[I�bY!�����{b8c>���m������l*����qnX-�b�ʄ����g$N,.�r��?�������Q9ZRq�̋���VP�4�Na$�<�x��Anܯ��{��b{�_<������������C�㈓.��'���!]@��8_���AE�6y�]b�2���@�]=���#�V�Wmߏ��4����o\R���/ڠ<���a_��r��W��4��H?5!��1i\�'�u�3Q��kw%��W�A������E#w�PY"A]���c�7�t[,����������I�l���F���UQ	��M����kU㹳4�g�ʆ�Sj�R�SU�e]<�E���_y%e�C����oU���YB`���hrv
�n�~��=$kn)YI=�n��V~��V��!Ȁ�SEkU���Y]Yͨ>eoD�gu�@�Ot�qSآ�;PQ�է.6%C�V�J�ͪx$u��ִM��h\Q�<������	��ÚDw��q,�=�?8s5�ȁL���ƟB�E��|�f��J5��Tٜ{��)j�iN�!.�>r�n�՛�G�/���T�=��X�{�rp�!�]�m��h�ݠ\�[6`F4�|�����R#��b�q���L%���+�e7�
�o�~����_޾ny�>��w�����/�!�۩rA����j�؂�S���ūX#
5l]����FE$�ﰗ�O�[�ϻ2��CPT{��3�ͱ�J�X���o�X͉���f�,{e+����|���+�#]V�,���KN0��x95�����r+E�#*.�C�]9,���%�J��<&�,�5��oS��¹o,Z��D�s1�Sk����0����u�����q��6}X�"�T@}�lM��� <8X�N��܍�Y���6��ty3陮�;��%�t�~�MKj�K�+�T������s���^�����"�
N���0�7Lo]�u����*�x�"s�U~�.������S�	<�%�{�+652�+z7[�gd,B��-�x���?������O����󽐃�W\�������͘�Q&b����%Yb����\`.aD�ek�d����zy}7o4�WV�/|�yx*�mҋ\<�]�}/E'��|�?��xÑ�8���,+38jk�xRY��P/���z���;�jH�Q�ÐjS�R�ĳ�[��Uذ�)2F�H~�W[g��B�B%b'�7�$78�& /F��́���sG�
��oNFrE@��mŸP��
��TkpY&i-YT*��|?���Q�<�_��jדqNQ[D�X*M!¢�Vh[5~��������r�Π����-/�1[]�7����a\3���@�IVdS��[�&����,"�)�Kc[!�F������T�z-��������>����z~�`�$5�B�Z��4����SF�^K���W�\t��M�U>BM�QƦ2Y�Y�rG^O�����2�{���*O��H�*QR{9��pA���n�L����ZP,�ǵ���Mߌ�"ɺ�Q_�ZqΦ��������3xaK�B�"�|7���q�Hf��A0=?y,���Ŷ� i����T���'[��y���`s �P5R���M,2?��,U�7�$Hn����I�
(�ܳ�pZ�dJ�K:Mbl_怭t��E���<7���y���{�$̧��N~H��/����!-�N�-yp1��W��7��8(���ĸ�[�����D�����Z~v>/~X&-��1��7�W{#Zo���h�<:)h��H��4j~��	� �
�l�v��}K�	�����39f�"O;�d�6���')|4�X9��#V!�I�,�/�M1j��$A�zQQ�	��IR�c�'!U�K��HB�)�#�/��ـV���w�m�Y�Bn�O��VĿ{�O�%B���(�=���$SZNn#
�s��>�)��@ޙ�5/�!Do�ÏHO��@�r�Q�����Q�{�j
Z%�&ޏ�.J[�zoD�����jm=㭅^̽\�6L�:��#����\��v �g#� ���+*�R�([I���ɸ��u���V�M	1,U� p�vfae09kK��+��*�6,��9�K�v�8h�G��@�<�2�hw�0�i�B
�N�m��Fs5@9_Y��G,/Ȝ���O��t��;ii��ZZ�D]�|��G�tK(�F�p�;�@�/��|�J�q^zy>[0Om�m�v�o)�����^�q�v���e_���/�����n{����O�L�����չ��(�w�ft�}���ٳ{��[���n��v��~~
8�+��Qu��7���/"�M��t�&?�Mp�n�[ٌC�@�-�0��(��uu�.�Լ�ͬ23���$M�;d�g(뚨�gU|�R3�_�)�?+��I���'A�������Ŭhx��6��%�� �!_�M��P*,�{��i��@r�j��j��xB�o�x���O��Ծo�<}�7}�T��� GC+�����.]9d��O���륭�ꑳ���5B�)�^$��X~Ҍ�meb�o?B��)�a dv��#ky��"y���m!`U�y�ve�C�?;�5������Y)(p�����/3���,W+��AY%��&�JЪ�ǜ����6��p	�ӑ��c�bk��H��d��	:�kVS����^+�� ���[ySmr4E������m�J�[���i	U~^���qk���c���?�q��C����J��'�%X��Z]��ɨ������@����qv:J����p,�ėR=E=P�΀�)4�-��?���K4�� �WȔ����˙d�P~�����:oX�7|���]�[�Y���}p�S��aF�[�[�F�������EL��c��t/gx�j�/G­/�(f'��2�b���De��1�X*e>���k��M1Z	��8��Ƙ���	�t�&4G�=cv�x9���@��A�T>�$)M�H������$,��0j � *W��f\��+L����t׉�V�#8��ԂI��[u�_��㈜��h��b����m���J#Y�sb��%���O�F5ӵ�iP�	�=�i��*|:u�ޖ�~��ى�_И)G�;��0�����@�䟚P��ތ�:|��ۣ~dJ���i�E�Va�Å�Ƽ_�B��,�!
�P����_��79&����ZZ��WFИw��T��e�G�qX�"ˬ@�z�>�ؒG� 1VL���p�2,}��L��??=��j���`a�W�-��o��E�7Ю���ݏ,�<�R��`;�,�'�D�M���־����)�fRO;����06����^�y�ˤ�=ϝ��XåO@��k��ps|��E�L�D����guO>5�	�ì��M�G�����4'��w�y�{/R��gkgҘ6�Ƽ7��Ҝ[�v�<`K���<�COT���:���ɔ�g��s)�_��|��m4.�p��+�[��Y�櫔E������P���Xg�o6�=��9�pa�����H�ڷ�K
�-%/�Vi^��u���[��"
�ZQ0 �g��y�9j�SiyfD�����qk��b��R�}C�8���+4 ���j��ߡ�>F���ܪ��ڏbm�zf�]��n�d�}�U�����D�\B�f�����f3��/���F@�Rp�Yz�{B
��5�������~n�&�l�^om1J.-C�c��\�w������ �-��,u�:��M2��P��@��ǥ��4��G�Qn��>�[z%�[����o2չ��>m8�	�S(�O�������[�ԫ���E��9W�ڄ8q�0�#���X򒨚B�0E�
�Ѯ�����7C���0P�pY�P������!�(�X�O���}S�a����t���?���������J7dq5�6Y�5���M����	�����Z���G�+\�w����:E�&~��"#n�P�������!U5�S�I�u����A��Q&�1��)�#Q��C����l�x٩-���|��P����^,������ྠi��K<�i?=Wɬ<1~�����ToW�7t,C�V�H����yD��SLX�J�F�Hn\B����簐�i���Y!9��7jרV 1���� ߘ��W�XT���$��x�$z���S��R7�"�H��z�Ԫ���cYrUQ�%S�0H�4��v�#dtʝ���J���� � ��߈�K&���^U8����ki�坘A�~l̷/#��K	���}���_9��E��;	��k>��-�'Q��e?���e���6��^���%�J4�y��,5ya�H"�.O7S�b/"�Z�`H ��	g��;H �NK�V}�U�TE��85��w?7gt�EOG#i8�'�"�V՜)n��a�x��ɾc%A�l��0��W}�v$=���*����� �zn�k�Oh��*�jW�݋�ix~c4�%|�>v� �М���F�*q�i�/{��K̳ϰ^�~?�G��g��qyS��A)$썖���n��h�rl�1l�ؾ~��ʿg3DH�W�ζ6ｨ$@���2I��}Lp�rvR��Y�����_�Tڌ���k)?���	T�����#��ʖ�R*���խ�,���;ޱ�&���E��^��m��G���d��Bq��I3��_���I�B��[�8��(��9��KV��4�uV5"��;�MD���q�9����ӵ�C�{�u���T{��M7���f�����9M��8mo١&��q��Q��Y� z0���X�m�Qu�Zɍ�B0�lnM���ĴOB{�IT2D�)u��U��*��T��2ԭ`�T/k�TAQ�^��IW6f��.f&1�K؅o+\��FNJJrG������m�.B�i�vA���MO�Lײ~MÀ�+����1���=�[-�yC�y'�f� ��)�Ј�θ��xh�ͪ6,��;�u�I�O�����*�)�L�P�~C����J����늻���3ظ��0���ZY���|K��t�y�%��"͆�3�>Rdg�3p�:�7��q":�@]Ք^Ь�\R��!���ف��Ķ���h}�e��ϟ��S^��^w�L^����B#�!��+��`�J�S�t�D����.��Z��,������1��E��@tڮ����B��:}K辅ك�'7ׁ-�`e;/�>�*�%](���U��=�Į�?��.%=?8�HTd�h.I�+��΀d<�x��`�� ��R\!{z���K*9�m
n�l.��2QE�Fg#���{����vH#�ڿ��>H�{=��L��02*�Dd_�:z-��n�S�Te��oT"����8!^����~7Z��`r��T:O�8�j�F�=X�0�����gg���u3��>\\ZUo(�j��������s���u���SP)�R/ E�Rʺ�-'?�@��ŸOY^76�����ӳ&X�x	�N��(��>���"���y�P�ވ�D<������W���6�������p�̳H��
�lC����j�1^�404�}g�xĝc�>��z_^�-���k��GDdɘ]y
��Wh�e����_�*���E3ڕn��w�L��#B^��*������@t�EH�/ˀ�
^���U�o�*`;Ӭƫ��Ҩ�:�vE�W<��䶏^T���O�{���Gm;�~m���ۭ	0�{�/<���j�L���YTJjYĈ��N��I��K�k�WK�>U���6�i���EW�`��K)3�t�}���p�g`U� >�ڮ	C�:�|�F�_���>��^��p�W!�����qE���\q�:� �5�@O�$�)r2�w *�Jپ� Yp��YV�a�$&\=1�s�|Q޳_B��b4@��t�� �N-/V�zv��=�7`�':8s�^�}���0�S�HB%�pD�t\��Q-�t�ǀ�Sغ�Z>�vr@`���I��;��hϬ�ؑ�'VH){�6�}V�yVy���2��%J,>E�Uh���|�a#�*E2Ϻ���e~AuI/wr�\	�y� \�Z������g����^>1-��O�E����|K肁6��7���2�h��N[�KJ<��dZ��W���§E�@O"�rE��<�fA6�;b��Ա  �*7�����Q9�N���&A��kY!�P\�K~;p�H�p��'�__�|�����΁�F�(�#"6Ks�ԃ�.KH`(�5��%A����e-���{�4�d���x_��ϴr�4<��tX㯡f�%S��a����~����.����f�q�������b�����M^�Iai㰁��aA�4�����W:�;��kn{��R�V�~�Uw���ޤ�%s�]��1pC������K@ѵ�[��4t�S��XS^N��YSc3��PMO�w��b�nY�M%K���pٺZ�|̗d����6m~J�-�)oE_G��S�k�	TҺ��k���2�Iyܩ6�c���f�o�!a�x��s�!k�P�1��~���p�m�r��i��D������-ߒ����s7hF��m`���:����>�?I�����Nۅ��F`��0H(H~"��x�4��L�zZ.2�?�j��� �q,ҽ��$4lI�$*��&K����c�9�G�����c}����yq���T�-�:=J!�HK�䕇Q&�3�p����PK�Ht��B��q��R���s�V�N���Y�.'�)l��S$e��f��v��޺d�W�3��k2��Y�+돆�����y���:��v�^%����&��,�-��r[<O��^��Vp
�-(q����m��bSu��D���a��b��wKB�w��4{�����ra�H�U�H���3tEs�s���C��1��_�������	rx����qs�Q�T(�d}I)犦RP�ӱ�X���@ȡA$�%���,1�L��q��J����F.��ɭ�=���h��� ��z�{'��Q')%N8^���������[�J^f1�v��J�iV���n�� �ȹcC�VE�T����geiQaW�f-�����/r�(��.��ރ��&�Z�z�a
K(����3Ya��=T��'��8�$��!D�[&��Ex�����	u�%�|�U#��Ջ�+ES��^�����d]#_3Ud�R�6<����d�]�7#��0��7 r�\ἳ����2z���ϊ����%K�(i� <��W���_�L�
���,3��p9o���)�ƫ$�PB`^++����.QI�b�U��6��Z�bԨ�2x?��Vi���J���}���PUB�+ڈV��4�-�,'{W����ae<Rt;M��F�A�KF��C�����R�M8`�J`(W=���rܧ�����F�@�<��E�~W���,$��!��c���B7��\�׍
�U�&�y����R�(�H5�r����6Zi���=��G�B=YU�0N�&՚����'ȴ�����š��RǊt�h�}�t��<Qd��/�f�q�4S�
���m:쏄��ɓ^S����ل���֤�5���R�������=1̞�ĳ�l1�@D�e4f�����O��A!�v�����jT�|��.�.l�����+6�!ڍ0�V�{�5:�{�Q0�
�c w�,"k�S���� ɡqI��h���yk��رTy3�o��a��L��No�����9w��-�E�%�;l�F���@;�{@W=��U�ו�����r�{����Md���Q��e
�l�h�9q6��\D<z�R0�]����Tҭ�g�)}�An��!�NRP�6r�p*�7q�e&q�1�6���ժh�.d��:9�����vaO�ꑻ������s�t��)�Hr��H��%��xѭ��S����� ��ەO��^��<��"|%G_�.�@c��~\z�,�;��<�6l@�;�iKE�'q�ي�v54����yB�s(Ce��>�U�+��iuotf9�V�]�K��>�5F�$^������x�@��P�GF���e�)�V���˹m�O|%2"�NN��*>}5��i +�8j;5q���w����d���b?��|�cNVa0k�%��o@����:d �f]čS��j�$}��9�Z�Ts,c�G����ހS~D����?�|LJ�haD��n��@��-���4��H�>�M��I��)RV�f8�2��&��ݡ�h60+ˋ����ЍQ�Xq�β���)Y谏m_~�����w�;���c�1Ư��~�RG��[L��H��,�m٢��d/�7���WL�/�Z������U�r�ܛNp�G1Q����2�5cy�~�Ա�m����k	`�n�� K�3�J�`��N��L�n�7G׀��Y�M?��Ft5V�Ѿ"�Pv��ތ�<(6^���"�gPj�aڝ�=I_���fV V�������[����W�������U~��73\z���M����ի٭
L�Z=��8qVB�,&Z���i����7L#�0�㩰�,��V��u���~���2��}a��C�\R}��u��$�	g��*����%��-uT�A�E�f��<Y�/�N�<5VS��]׹�J������EK��n�@�f�����P$���\���`9St��tes�g���5���{G�������z�|�ke[����ߞ�9ķ7����U�M�n�[T����/eTō�����}
)z���p2��>uH V���	p6<-vɇi�q-[� RS� �09�EϺ���)vE��k#�E���S	���kԡ[Q����|�Ջ�V�2u������e��TNƂ|ۓؠ<���G��IFs�x4��JW�L�XmK���ޟ��x��M�J�_�1� �h��u�Y=f��+S/�8�����d�0�t�� �N�Ճ�Aw¶��$��yݡG	����[�p��i��gA�{�i$�,�h@7�r�g�N�ݍ8�3��K������*�iay�Cl���M�2�)����EOԻU�|��&D�5���10���%M�F��<d������W�^� j���Q��D?��:��5��+�v�|��{p	��Bh��}G�Ȁ g6`�nM��%1e��4�:�M��>�*(���#[y���TMc���sv3�<���*Y��O=��Iz��U�Q'ճ�Q"�G�$��/N�:k?��9��86�4����kG�ٺ`,Y�a8n�a��j�z����%�E��|��0�����d�Ǧ>'�>>�&;��q�2`D�?R��n�0��� 9��V�3i^��W��|�$S'r���2 �B�A��y�k����@ȸ�KIFƀ*�cQ�4B-�E���o�<@@*c7�H"��T�;���.��|s��&��tͮ��(2�-�O������G��w4�M{�y�!��ua��p����)m�aS� �Re�'�� ��t>w'������\�m ����*�0t�K�	>\r8?4����b�sh�w$�n�����q�Ԑ��ܚ�gLF쫺@�c�Q�7��6cR��Tu�&%�5Pw�����ݕBg�3�kj�ո�����J���k-��	?�.��0���
8ϏB(�F̚�`�e�0C���L:B�TB�Y/�����S�/��[��Մ�of���xG�|V�h�D���KyA6�6\f�٩��/P�q=n��o�|�yꦺ�gr�ak�W�����Ee�q?���񔦩�tn�!=���j�������Ф��{�=g���rSj��P2uvx��T��/4���MXu��L\Cy@�?:΀=������|9�(7�����D,�� йqu�ů�=`v�h����� /�i/|ƪ%J�:��-=�0�"ɋ!��pf��i���u�B���/�� �^�[.�2�O?3���Y�>A��C")ۑ�{�0$maSY=�����ф`�"�
�Ħ���U���ݭ��2åws	i0�'x����T#�S��4nY+G�&�'/!����	��Z�^�������3�58K��Aj�y�X`�As�+!L6�����4�P�~�� S�\��a^�M�a?�h#Pllvc2� F:!��.�f���d�$�ţǥ�/�E�Ey� �f�oC�������Gr�j�ƀ(mb�YU�c�q=r~��-&g�Q��n��h���ڿ�l�~y���a�S�����|�/pI�S>�$���>�� P�>���ұyc	�B�܉���2(�(���5X�2��OKS��޳䆮�a���ف��t�oe�)靽�p�No��O[��y��u��&rZ�#g؃j�f�=7��� (��4�(�31 &�ۋ�eĝE!K�	��6Ȣ ��T�������T뒷��#)�G�d���|q�b�����:72^>�>�$�=��\�<8��S,g� 1\�8�J�<���Qz�)�^��ɣ�Y��f�BZd����)�.��7C$K7p�w$�*��j�<�-6F��0��^��̿�~������zTG��n�+1҈c�ƥ����~�7�̠o2�>�Zr,��^>�~�3t��ig�:i( �aQߚ�Gb�p���=�.�,�w�,䐛&�}c���L� ÝR��c�x�2r��Q>_ªm�a&�;2�(��a�ӕH�q����K��z.ؤ2� ��=j8�]��p	�:�l0R���?k����Ð&�,<W�M�z�Sѷ*�����m��]���J�\>�8�ӭw���X]mW\���_a��f��$���tӊ6ԑ^����e���@]rMO�$4��;+�zs=X=�&�/DݶN9���J43,�w	�T���E��+��#�>������9g�� wIr/�+�B6���{zS"�(��FH[���ea�Ŭ��F���}�s<6�o�`��R�ڸ�I���<���y�Vu��$�<�k�W��A�|ft�N|7/� o'�τ"FB�q2�y�i=|਀�i����+���S�����&x���$��w�f��aCa�M�2,C�k>q˚#����E�����W�U�����?G���.����g��|:靃W��~ ���g�9�U�v�a�y,?�X�/�ⱞ˶e�D�՚j�s9RY�V2�(�:�=�~H�k!��EY�˻�7#"��F+�(8Q�#?`���;��x��+$��fI�Go[�L@kl���ԈŻ,��z�|K���N�{��ni�r5 �(��|�!c���w���.��Q^v�!Dd^��U3����x%�������A\��|�A8�]��g��fet�O �N��Uξۧ��"wru$(�3�E���.`��t٭HΠ�븲Pr�����:�hh^]>�����j����N.��q7���I��6�g��Zp�/�悩����"p{MDL��mW\���S�`���C��BmEnpE.�d,3N_X(X椗uYρ]P��I�,�Ǳ0|z����pHF��XIKl�uj�?l^Ȁ�0+}rF.�j�߹��T`woQ9auW��$\��W����������_�P�x�����hEE߬v��Q�j��B�����K^Xyl�Ɣ?W�Wˇ[<Kg�r��ڋ���dÒ��.��1ƶ�۾}X���
�q��, �J~{8\JV��Gx�q�OE��@�.+�zL�9C��{t8#ԝ�����X��'��=K��(FĲ#�7Xd�ǝ����@�� F��V��gŜ���2��#M�"f�=M�z`��ff�qK%\𔛂�C}�{�본v�F���������S����z�D����>����s\���R:�)����l��Uփ����Y��lޛ���}����j�|&F��7K�4G�<��H/��c�C��iޕ�ov�V,r�b���ՠ}P�"��ml����/ƍ1ʤ	� p���At��o�RoP��]m@��4j��*��q'��=b3h1�4k���tg�6��;��l��3⎭0�Ќ�bN��>���.�vF�
<'4���+���rBW?\B+6��ⓩ��Ӆ�l�tLnN��v	�d�����=��,F�p<a=/T������U4���So��7��d_Ɲ��d�sm?x�7i(�#3y�* Rr ����B�$���YeWI�ѾWS���Xd�"dE�`.�G"�e-��#Y�)�;��L�l�����M�
��62Sx�l��8yЛǇ��IFV�1LTW�	%�����3t3���Ԁ�^9Aܸ+�:[=aq[0O:�O�lL)��~$��?���#�����[Z��=T�����*��;�y��`+y��DQ ���Mr�{3e�딆���Yí��rÎ.%j�@��0��?"�8�R�@	���0\c��ĩ�q�h���,[��~����Ի-ǳ�����7<���5i�����}`����
{uۿD��d��I��lϖ� ��cq��\w׉XEZ�R��	 Ρ�޴�C��ZB�_=:�չ�U��h��(��㘿=LT�d5w�c�_w�ׯ�o98z {z_E�֤��x3����f��0_I������F��W�rB����y8t1���`�8��~('v8V���ȥ	Q�2n��j��//{�>��$^��1�4Q�+|�]D���ф)W��8�]mB�9�l�*�j}'05h��� ̷sk�;!�c�z��c����J��|cn��x-6�/~�Ƅ�y�c5̀���x�Zj��R/�^Put�&�SSD�z)p�G�>M��1��v5��`����1F>�{�������+��n?pH��%�\$^�{��J��~�x���馟"�<��2H�����=�wV�򴀎ޢ"u���Rڌ�j�;|.}õ�ݟˌ�",��/碡!��:��K�P؄CAf����(��KQL�ل=c{�����S�75��{�:�����=���pO"R`�}J�i��+�,��ވQ��k�s���D�5������.8D-:�s��2�HhCGc�»�u�!��m �c�� ��J�	�`��fa�w5
Ȯ1��'��D���q"A�#4��G�UĐjZ���V�b>�2�a��$��8L�ZcQ�C�ɩ1|`A�����좕�z��]��:��ǳqm��p�LIoU� \0�AX�>���K��XMA���Ǒ,����x�����K�e��,�aM���ҥ�ta:�'���e��Pj�IA��~�xGX�F�וg(�8<�q�p�gͅ�aﳒ��:�g�b���G@n5#]c鲵V<�a�Z��|�Ъ9�U��P�Y4P�ي�#9���f�x3�݉[��7zW�V-wU�&"��ĉ����n��t�Pa�=ZE��Q���Q"��ǭ��[�r�)��m �A��W�?ܸ6�Iv.%���%҅\����~$�3��������?Õ�N�k�� x���pfx��}���W(,�	4��\��E��x�@#ꚁ�s#����'L���LKm�P3��J�z�r\�/`������4`;��e�\R�Ί��s�Ͼ!��ݼ�oߺ�XX��3�����.��)_j��W���q�%=���TY3O9tz��#��t��b(^��w�ݽA�'��|�����=CՋ���a�#�]�4q�ɻX��풩��Q�@yʠ��}�:��C�N9)���?2��I���O۩'L�$,�X����_�
�A��?��e��>�^ڷ�`�)��JR�l3��v�O)2Q�kC��äf�{'�nAp�����L�� ��"�שׂ:!6tؒ��������S)m�v�-�w|J'��]��B߸����@�l�<eID����v��͙��a�&*_פ�v��v���~���R�'�"�!����T3N���S2馔������5_v��^9R�k�����/��c�� ������ݟ]�Mmu�p�{�iG��_������𩝪����wur�y�_MM����vu΄tBP.S�	��z��w��E>��RzS|T���MN�AmqV�A70/�����:��]3aE� ϓ3����N�q�U����q ���+�|)��y�ke�|��5;ZW��˔\fWL��Z�������cUJvv���2��3X2le�-^2+� _܃9�To�y��>a��b�9C�P�0(鹚FM�0��Դ�x;�dL���Aj� �9�����7�^$z,@���R���&ŪY:�8v�S��-T���~������s��M�g�R��xw�J"�8H�C"<��T]c<��n��{A-����C��S3��M�<����rt��mx�.�ES�����7����I�eF��i��Z�i��,�"��C����c^�802�x���� �?����
+�"ւ;@�,m�\�[(;\�_D���C"Y�ib���LnR�}���|*'A�)�o΂���qt�2t~(���� �D�����Ԙ��=���\dV �c�Ig)#GA@1��xp���uc>��yݣj��m�5���V��g�|�%�tE�ktnf9 �R��W�.�K�+lE����<?���Ǹ��*	��{@[�S��X�۽�bL��C��S�-��!�Od�erH�4.;N�1���D�A�sg. ~��t?sL-�
D1s���:�=Qj6�Y@59zUГg*%���@�*>JT2�}4�}���+����4a�ߪ���	^�W�?�˜c��:�X�ctۢ�k�G�UnsYu��j	����hӿD$F 
��b=��95�����1`�9�f��=�&FA�K��y��R���G&�+䔏�#1�G[+P�����%�b�C�ʴ~�<���E�
K.�n�L ��Z�|�������d=�����`ET���oU�έ*�T��Nd�*�}�uFh��`N8�~�~��:g=>y�Z���Հy����cK#�=�ūRGD��@�� gu��&�R�_{bk-���f�0gE�M����w{��s�ΪA��Ĩ6�|�)�ԯ��'�
>N�"�e&�,U�܋I�.p�T�Wm�I<\:US��hi?������� ���ү��8S�,���0�����
Y�����@䒪�_e�ЙӃY�r���}M��%���m���Dq�1*8͋NٻY��D6�q1Iuf�-:�P�Ć�49z�=�$�9�ca�+M�U���Z;-4�w��1����u{�����^y�c���7m�S�����\��UG��[������SB�M�EDP�iF�[���9�4�]{]�m���c�uP���;op8�[��;;�+ZxB������i�ډ/��0����~���U��^Ѥ�����p��N�Z�CЀ��g���^,�֕?d�H��R��	���!qV����2�S��>��5�\ȍ�{��p�x��<_�-C�؂�"B�_������9���;�h�v�un�p'1%Y����O?�sڷ'�i!�\A��=?0S~x 1���Ѐ���D׺�,*����߯���^�Z�SR�&�;��i?�L��_!9�.0��z�| Ig���>т��3Q�(k+N�ݑ�\��9�ʢ���v?��h0� ��d��n��":�6�I�C� �ž��Y_��"������.-�8)�(Z��rq�,�1ش�@T�����_�~1V/rj�aB%T�X-���.��4��6ڧ�@��V�2~ �ɝL�?�/��hQ���D�6�(Y��P0 �M;��fǬ���`�xj�oc	K��dPd0l&%G�E�h|�ŝ��^d��3�TI�	�ˉ��1T�O$�!�)\��=���}���<$W��7oEDOS5�;C��u8��+'Gh\)�压��~<�Y�����1�#�n�(o�]f�F��C'��"�p#z���(��-3���R����Oʫ�1R���R.���}������b:a� ����
t��j���B!��v�|�d�2��w-���m�s�D�{�`P�T����i��V{m����u00�kX�<x�M�R_J��Ό�� ڭ�6��=<:���$�:}��������O�U9�]%/+Z+��9�/Xb��G��9pV��G���@�*������F�г����i �h��0�����i��*�2���%��1x;EL�wM�K�cx�Pp0���#�g_�
��Gza����l^�YI�vb�����h��������"�q����[aC<ګC��N��MC���^�� �Ge��kq����E��r�uƝ�-�����1��V�u���T�5��mڋ��n*���i*�~�E��i}����4,<�I^�	�g�R�xZ
�F+i-�#Vy!�[��u��:XF�t�7\a�� }^)b���ڔ��FE#���nt�0�HH p/���<�I�4�+
7/�
�.������['�f�+�O��$hۻ��G�K(R�F#AL��Kк�e�����B*gD�~�x��&����h���!����R���zf~en;�������1����~����pq�x�
�_oTP몘g{̿�\m ry�Ÿ���~����;w���������_��t����~���M!>�t�:�#ň�6���Ź��d�ZL����k���`�OL�UŰ�:��kT#�[����ǃ���_Zv��͈�����sK;ͽ����ӹ�({���<\�z-#���I�˶eG)m��b)`��y[������`��@oh�.'��u�a(A����g�q�!�f���G�����`����"$��Xe��?��yi���<����5�2�Æ�o-j�w�ԭ;�:!�����Y�qk�-`DV{ɢ@͊ h	�W�,�qF��؜t�BB�N�ylN��'�[F]�+P�3���b�W���_�P����l���PDK���� 4ܘO��֓T-�c7�P�룬 vp�M��|RCIA"���o���8�Os����9�����5k�M�Z�4e�{��f�>����C *�y% ��ZS�ʆ񙏻1p���Y���/�����Ɓ�9��Z�X;Y8��ӏ�g��j��eC��p5�AoR):W���N���@��k�2C���<���H�a>����!*��ث�'�-�	/Ij��{"�������?�x��9����#ǢP�!���u�c}�
��+yqvL����N��=��]$$%L�C���z��N�<Z���E��c��.h�S�
�c*ɼT�/��\�@�%-!��Uk��M���`T�T�h[��ȃ����:�����uf�u�h��<:�*:/ѕ�3�8$����
��o�$��'��o�HML�z�mX��f	�����E%(��󞄃�Mݓ �t�`�����X��n`�9���gA�K8��M��fl%��B|��:��ȷ�4R.�-�9�S��HO���C7��TDt,���W�8����3Z�k���]]纚>Τ�b!��b���Bwu����<&F��/����b-!�9$��u ~��tI-� ����f�K�CA�y7Tl��O�6�[2w�ӫ/
Jyl.�"=q/`�(���L��kAz-�a�|��xJɤk���#�c[��n,��,s��ȍ+5��{I�ԅHPk�=F`��6��o���+����g��R� �i{�|�]tZ��m����	��Vs���u�|�[�vi�0��6�����t�d��Q�?��'���E>��|xv�b`��Pv��]E9��A��vM�,*o~!Z ����w;�h2o��$t�'�$��ω�hC���ex
vc5���T��=��I��<�v�.Ɖ֮�r�hl����v(w&(�b�l9j��H9��Is7Mq̰�.)!SE�X.��gA�u�Hr��*
���k�)ź�������eǻ�,Y9�v�q�"�V��n��ԼAg651��q.���h�s�=��ɫ�f3"�^�:�y���	�����h��@k�e�F�����f�ӛj�y(�Iā�L����(՜�1�������d�ӆW.}�SS�'h�^e�o�ޑ������0��_����ӥ)�+"(5+Fi|	�q�sΧ'�����������yd*��琍�A����jC��O�D#�M�8&�;�$k�1OS���P�j����I�࡫���!�t������zo>=h!����;��W��`;�a�D6� ���l��������Oܼ�\n�R�o^o��Q�R������n�C�_�c�n��ov�\Aư�c��s'�%K�D?�??2���s�����hn�<��8(��,Bʾ��e��F�Bsd\�z�,�ʎ���
M@wI}n1�A�k����ѝ�<�@g�`�PP���Z��;��Ll�i�<g��Wk]���ԓ&D��Y/�t�@��y�]�8�Ns5��m:;�
���<����w�'��0���[��Bd}u�tLZ��
�*������{����vA�d��v��uDi����'��&E]�L���x���_�T����j����0�3P���C-)����aK$"�~9�R�f~>aFh�_�9V߼����uL��u�e���P����	�/*|�.�b�R����x�a=5@�K{�A�>��:*A�tI�u���{��p粣�,��7��ٍ,<+'�-@5[�'`���3Mk���{��1l�=�e�R��bК>O /v�x�m�̩�3��|G�?�����$
N�yc1"�a��� ��vR��%	[ /���>]���郎a��t�T�&i���)n<��3H�V�o0���/���M�`FF,����\��!i>���!�+�z[��&�U��]EHM��4��1���j���J0�.�:'�wk����/j�����'F�\1|0�zOf�#��~���Xև;!a]g`�B��{�V��o�Ϻ�p����d�y��+�46��M����G��G�v��QҚ�z gN"�)�{^W?{�@^^}�k C���@u�3���_����h$A��7��Q��f1MY���Ķ�?8lJ��P�
Q�;Z(������8��`��5>D��(��2��E_�u�4L9T>[��ᥫ�?�tr��,g����F�鹎�E9U.�{/������}eR����B+�����N~�I!>�r�b���Q�n �lG�ص��S�ׇ���A������3Y*b��6�L_|�M����,������ld7�im����,���O�m��w���<�[��n��ċu�U;t���R�c#��Vo�W��6뿛��Fu��tYe��q�A5Q������!EM�
����/{: 4���M�#?��W�lZ�ɇ"���&9��v�ҷ3v �Ck�Q��3��D{�� w��&�8FM��O��J�/�R�֠K��춻M��4e~�|X/�*R�ѹ��uK~`�*_8\,z	[�#�)��Su+	VA��n�ڒt��M��,��.2�?�0Ŝ��UwW7����m�̀�	���n56g���\�^S�ҳ�~C�%�BWv�5�U�H�"���ֈ����'�X����O�PpR�����xjr�(�4��9�*c�|+
�;�.sY�4p���Y���Dd�������b�4뺋������W�d��
j���!A�����-[��&���E�����"���x5G��U�X�&�6
鐼@�7A���$��O�.l� x��
D
�HY�w�o��b�.�>Y�Yl�
h�>���3?�,8~Z}c�s)��^4��d�)��sm���l #i����q����c����
�mұC��ׇ)�I�|˽��['�&�:�1��p�Ҁ])��#)	.mI�^��z���ٯ���BZS/d�K�D4��m���EQ`���K`��s��k� ��n�����G"�W�W\���ޥ�I{	EeNa�*�-��׵Ha|sY�����7ߨ� -�R�Z�4���;"U*p����G���J�+C�����{m�BA���A�ܖ�Yq����y��+y!�	���d�Q��Sf���x��쾎�-MD^�Y�v3��P8�49���,��Z�dq��=s5���|=��b!��C�u�uV4�OgY�'��z�!���NJl�$���ѹ>D��
�ls.7߷U,���T5�ۍr��s��E��"��lR�u��Z��Wy����m"b=�v�Lg�0��}�V�����<�+8͒�+mp��k�Yq��em�E�/V �.v����� ��4�:�$	Ux��-��#���B���dӴ~A��j�i�T�3��pmc�RL�`��"����+�8�4��T�����OL��nCCNb�z63�$��]k]|�Ӽ,��zL��	MqW���7�(�����T�co��D�=J���}�plk5Uh���je�ˑ�jK�.PѽM΂PZ�{'	�������]�IN���?�ud|έ_���8%\���%*�����4-0��P����uV������f���}��~؏���[��Ƒ7����)��Nɏ�v�x����b��$"�Z'�IhU����T�>��i[`f1ɠ����V�3��H\�Ϡrd-�5���1+�8DMQK�K��b��H�О��[�m�DQ����;��`�%f�nA{�#!txI�OR$G&��L
�Z�5�ھf$Q�f��IW�T�����t��*�G" �X̧6V�o�Հ���� yRR?�������Q�_�J4i�����x_�e� ƭ`2`� �h[�;������ɍ�&�Ϭ���0��aֈ�f�;H��"�uI�0F?q�Ԭ= n! Y�A
���곸I�q��kK�%t��!ɬ� a�լؕ���0�A�Liû�Y��ɯ����s���j�����R��f�$k|	��.fW�g�\�,"�[P.�����f-�Eh�Mg��J|�*B���7;�l�m�:�;5������������6M}(��t��/��?��߈� #��e���&,�'��.3�ZISM�_�ϓ`���KZ�O�����N������KA�;VA����(]Vnq�l1�����{	 aY�=�j�wx�f�Σ�Bm�����<��5����|�q�|��>*����T �S��/Ƣ�.��l	,�?�g�j5�@.͐q�tD����㱌���M�͟�����,��Ƶ�c�w}� ���-�/�"&Q^���v�L�I#�pp�	����4z��k>��{̃gPu����_ʪ�@�n�ϗ�j�F�\���Yɞ�:�>�z�2�|�:��F� b�A	z���ߖff9�uE"�EF�b������%BZ��M��������8.RH��=D�W�l��w	�<z�5{N�A^�*����