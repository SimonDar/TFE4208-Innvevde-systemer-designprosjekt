��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� f���o��ʽj�j��d ���b�����LMh�Ճ�i��RB�F~K�=����x�a�0�l[d�{�y� Whkܧ�(J�AS��x\T�Xy�������@�{Vq�ܞ�N���{���v��|��7����҃��b��Z�}|G�ܳ>�qC7�vv��h��Ș��r���h��88�O��ET�Q�o��WŐ)bB[&�B�(���U���8jVB��27046Qvr��]����tK&�D��(�������]�֊�.��H��J~V�zU�j�\�������#�W�^�y�)��k���q<��z�4 �.��ݧY�����{�$Î��L�\�	�~0�x+x�3�����'3X�L����
Gk��x;��ƺ'�b�z�\2G?�9��r�9��F��̏�Љ&pp-��[�hhQ�:P��{���U ��~��TAطV����]C|��ڀ�m� <�cYH�I�*�~F�+�4T5ǔ>��%̿3�ͥ�T�M>��a�h�J�~0�V6yv�1�;���+�����4�wbF����Rҕ	�3��]\
J�}W��Tm�r~��;��@���T�~���ߓc\�i��GD
����}���7.�?�Γ�T*�Ȓ
���O�� 8+����Z��t��|x!�s��k|Pl�T�]K-��h���xcڸ6�I����N�������JYid���_�<�ߊ��3&4f`�h�;Y��ARS�d�N\g�xw��_��]w�_����#Q&bf����4y�L�~����5����ZV��T��@�X�6o;�:�r�Zt��s��h;qL�:t�����2�D/��8e�9�\*��G/  ���c����Uq����ܝ?��繀j>�sà<��}�x�HJƒ�D�乼�wͮ��$Wǋҁ��z)�+�]<^���Ҿp�ui<mc���_����������2�͍�L����X�M��;|m�n�U{!&Z&,�Sش��,"Nh����/G��,��E\o���<��R6-�s�V�T��'a҅�c��ܽ�scA������<�_�N��:a蟻l[��m��z����^)�#���	���G�X��,�Z��F	<�� �cK\��1��Fb4�=��q�i�M���m�%Q�u���%V<��J���`��m}���iг	l�L�W��a�'��
�o8E���2T�*^v�k����V��������QL>�����\��p�v�R�O��1zI�GTCH�C�2�{2�Mh^�\F�@�e�wlh,nN��np���x9j?5�e�uq: �S�;�o2b�쉊Z��o�2�1|eE��� �wɗ<īa�7ҡ��-�y\\���������2����l��+J�%+NG��gU��5K��h�H��������x��-5�qu�٣��U�:���ܣ_�5���=�^�HL��F��D�q-b�%L��!�b�o��� �c��8��3*�/ˡ�a��pl�<u�:X���?�'��г�z���X�y,�S~9g[�7�Xɣ��0j�+��8�?=�mo� Sӷ:"� .�xpHҳFH�iyd`i���А?F�[�G9Ny�k��}��Le9�6�j���n�ဎ������#�4vk��LH��|յ�Ií�6=5��=���;�����9���Б>*؜`���Hǉ݁��?���R�1��FS�����Ͽ��	z,{�P���z�_��>�i,y�jy`lQ�/�Iju ��m��5��V���q$1�ؑ��]09<!~�miQ<�ȗT�k8K�B��'� 5�a._Y'N�܀��Z:(rK˼�} yϑj������F}mA��W8�
�����!��*�	<9�"�>�#���v�f�~�3B6����/�|���/�R�,�|��3q#wP�w��.o���{b
R��
��W�:���U�p���܇JN.�ݍ�
h8�]V�!�o�����w�7�;-ђ�z����ͯ�a̸�U�4F� A
x`��1���Ym���gE����">*�̘L��p�A�������@�s��,l�G ���]a�.\�Y403{��lq����P��mv:��͹YaŁ��N�&��|������5�D��4�l��g�Џ1=�x�C�1� �.<������Bv|�����g;��ޚ���sL���/Wvԟ��H-:U5ҷ��͕J$y��
��h=G�6A�Z���XӟZ���EAb�&��4,�{xp�"0|tP_HJ��:��F�ŷ ~��N|gt'�oj`,r���|����V�b_��㦴�'�Orٺ�!�z��>u�$�d�W��K��V�n�w:9��"��\�d�tT��kn8J^v�mhߚ�e�T���/�oe�	?�x�RMl�ڳ�m��B5��伥Y�;�$w�Ϗ�^J���Y͹����;� B�c[�!�k�'��˺L�tF~pE4Wy�ڸ����j?�Y��������v����.Ȳ�l9O.$r��7%k�#cĮq)^�M�nO
J��1��ڦI�,�A0�v|G���H6���h{A7��;�PYz�;U$�#9��*�ЖT��VV���br4+�B��kk��M������Xn����JJ6`�(�������P/�v+�I%�xS"�m�N�^���8K���i��ۥ׫����[Jku��8��]���p���������^�L��/�?E�-�嘳Q�R7PE6]E�l(��/Q��M��Nl��c�%�=y�-�'şJ	eT��P��e�=)�]�wDi�&�LM�I��a��P���h$�x�)�?�K��l��|�MS������۞�;�^����(K��.��2~�i�m#�O���=l	;��]p[��� ��<�����6�do��mE}ރ6�K�$�L�j+��75,�Ia�5����0٫���O��0|��L!�e�/ϔ�c	arU�@�$U��|J��<�#P�A��v�H^��gMz��]gٹH^�y�»�ɕ�L�#��;�Da(%}r��䉭��O}��jb�pѫNP��������s���LC"c�s��欚 ���/U��?^�ntV(�� oL�.��Umb0�6C$}%P���Fց��?������ A�I�ۡ�'b��h�E[�)�B���~B��0o�	ߥu�_w��ف6�XJ�N��l|{��	�l�SV���&�d?F2�^���d���K������Z	��'_��j���3��E���.�1
�}<K�{�,�.� t��(̾U��K�t>���Ըac�IK��\7����Sx�bs�f��E{B];�����Hz��ԨiW��|98�oh�{�ԏSf�E�Q����y�3z[7�"GF|$#���@��˭� 4]�T�&���������⸷�s�fDPς��0�`�$
��6����o��N�)�\M^��'\���rߒ�<|&�`�#�s댇����`�w$ *� �i[�Q̊?�9��?�6^�<��[Y4��F���~$�$G��<7ѱ_�d��!��M8%���茟�%�,L�a� �2�]N0l�����j)@H�HUE[������B�������P.8��£�)θ&zb�k�>5]��d4�_6�m#iG9�e<�	x�܊�/}!&Xǹ�Fi�N��Mee*g!�D�������FH��
"����_T��tkQ�Օ�`�~!��% ��цK\9΃���]{:�;Ntt,)���c�|���=�?�I� �[��$AS2�<��~�l��O,��	p~�W5$s
׫��b�yс&K��ܵ�R���s��z�U�
�1���s���E�3���m�(S��ΔB�N�I�i̠�P��Q�%���?��I��ޫB��ɠ��k43n}c%��?-a�a�}s#E#"���5�?5c��~���Tc�̛�Iր{k��R�2MW���ga��հ�ʹ}s�OV�0�1_�(2���xr}(W|��o,�1��aݐ�	+z%�(�v���S
-_��+��LN�;P:�4p%@����Ye��) ��S�x��	�n̿��!5�I���16T��If/��4�e@R!<{e�-c�bm�/G4�6�ψ��!���,�J�������*�h����Ǟk�j�.s�׬? �����'�����=_"�i�(�{{��o��Б�T�	(.o# ͂b�(���N[��_�DFV���u�PGS�v8��Q�&E��	_���S"w���z���W4�H?�'�=Oi���Um�K�Rm����-�X�=Ki���b�W;^#�>S�8�R�'���nJ">�L�i1J���p��-y�S^��������q��
�ۮ���"D��Q���z-�K�`-C;H����ϔЛƯa������X��1������.�
}�|���Ⱦ�Ցʥ�)�ũ�F��]u�H5*Y7ӟi'��]B�r���^1E#UV?E�PVJaͻ[AňtuS��aN/x5���-�Q��As��aג�s��U�{žᑗS#&�<�{�_��6%��5tUZ߹������ć��m4�y{s,��~�bS�"2V4�9o�l\����QiC%fLP�h5vy0��E���wx'�rl��-OPm�ʎ6!�� ���I&s ��HO�3*�+�2�K]��+#����ʟ�g�g[ZD;��ӎ�7,�v���n%��L�k���j�,�KqZ���A��-�J*���77�>n�������)�:WrD���\���x��#�Tw�I��L7 ��c|�����`��;j����q��B�c�7������p$�l�B$����� OO|)���8��aΒ���b���Ac_TSA'�_��Jg�{��q{�*= 9���r���);D���g�ŢL;�Z��O0:02�ld<�!�(Y���.�Ǫ�F�Azz��ҕ����9'���g�.�}�+0ov�?(����3#
���k�R�U��SN�n"��$�d�ԾM|��e�5��X�#7'��V`T�H����B��B�[N�A[�.N_DX�N�`};V.lM��7��Ge
Ƽ�����\�hlf�{Yx�镜/0������*�Z���P�lE �:��7f�ю?��rb�Ǉ�jtw7��]'�����^���E[�ϫz����x����m�8&���_ $�ЃF,��d�v�� �~���.���<vC�r�r�<��hv5��*��*��b_�-����@�>G�~0 ���cg%c�e��#��ǺQ4rhCؔ��vY:@�8,�PvTED�9��]:�r�Er�c�r�'����r	Nd�1��_���Q/x���"�~o�o�>������S90iHl�szȳ���A}�� .�q�p���Nt�g���R!bp�$��\��I)Y�f�sP�����\�n��A�f�lrtQ6�!1̐P�ĥ�u�H��.�[^�g��8s�f1�s���߃vʦ�+m�ܢ
�����p�tG����JL2hUB�X�q�3�q6�*F����
��D�0+���8�\+G�ȋk/�_l��IuC9����)����	?���|ʅ꘳oQ�] L,@̝N�'B�����d(!ø]b@���|�TD�h�V�柋i�9�1&�5,��捷��AG���D�6�v�e��L�ӓ��%CɊ�T(ܬT�EX����u�ʊ\��J��]�I@�J���E.����b&e�Ȣ��������X7���,�T|C�uu�[`[G�h�|P~&kSL儺��G�|:]Tہ�[�5<Os/Q�O>G��|�+��C�5��j"|��;�xU�5?t�
D/�1"v���L	�r�a{J<^�N/�$rQ�xN�J�:���Aʓ��E첎���6Ra�5_6�B�+��A�y��p��a%�Lsq<�����G��jj�܊��N�G���C}�q�J�|��9�L�}6v�����"�����Qp�5h���'�;?�Gb�a��R��*J79�}5����	 Q�-f��m�H�8��$��y]�.��>T_�O9r��[J�-"F�����}�2I|�w/*��� �n�o�x.���nޫ�_EŮһW�ڛ��}7�Wg�J�CR�bv�vU�����ƌ�Έ�j����Y�d���m�ܗ�9A�T���2]&�:��xc �)����%��s�$\�ŝ�ʡ���7O�AI�k�mА�N6d�1=aQ�T_EN��R�z��ʋ+8>�����`P^%Y
Ċ+<qI�9/ur5�`�{?��v�tc U����* ����ȭ�z=�
}_���s�99c�#
�b�hO8P��eՄ���<nM4��ͤ��H5����j�ӵ������%R@1���~D��|͐YS�`Իrp�FU��}��%�QGk��YT��d᲏��b����Jh¹R�6kZ�$�8��\��t�芣P�i��(u�C������_�Ų�a��� ?'����@v�	�~���W�[��XӅ��Aa���T)�A��Oː���S�}_vY=�-�ܖ�w_VEjI�.�7	�������n�,	�V�I(a�����%,�AC�Կl,Ѣ��ա�'d����@/�g����$1�X9���k����Դ���;6��L�r蝚J���ƶq?l,��E������*�ɿ�|�Ć���K0V���ɽ�ؗ'iX8e
�V
ѵ�"ȴp�����_t���PG�� aIkqzy��̏��Y*v�W��o(k�Z���t�-�9+��+�Qs�/�:@lC�{,G����vol�T��e\�D���l�<�H���|=�
�����&莘.r].�%V��e�+��:Ѹ/�3̼��$���&���/�*o������W8��Xg�x���[�͂�]��v����'w��7�tǇ{+�;�y�ŬW�,�q�x�8�d�	�n6F@��،M� �d��&�- �0H$����y�i�K����*���)h�z��CH��_���؋w��%�NW���zmί�&�Q�c���i�S^4Y�I��X�l<�y��;Y���T$4�6|��L���!���y����u@���� ��i��!<P��ں���k>W���ć�5�W"���R�t�y���=�ٻ�:��>��V!�4���-����*[���q�0<1����-�Xߒ�p�w�Z٦�(\�F�K���?��Gm�/��L� ,���R����jB����싋҅����U����͘m����}�i|MS$�j���2��c5���sD�u�j�T����OS$���2~��䝼{����B�`2ͅh�nΔ؍�C���c�xZ���(��d�ʒ����u�81�c }�0��X5i�[P��h�Э5/�a͌�J��2�g�ŵ��\d�F�}�B2�j��O&��vp�0yrJ�\�E!�/�!��+����yI� ���X����W�(���������
w:��k��BUSq#��,�������SJȥ�$���Dŭ�/�
i��i䍈*3c3�Z�'�=Kn����4��lo	��i��B�%���ω�%-�T�Ir�f>0�7*�"zy..�l���G%X���e���8�
��r��|/
�����$�q4V/L�ۭ�/�g	�O*�Ջa
%7�;�l�'C����{�gR�2���߳��*,�P���l�R?�~�Ӹ^7�����ޞa�ڌ�:�2��d����?��*
a�����Q}YL٠Y�߁_���!��"�^S��H���Ĩo$�_��G��"�Z��-������i��D��$��U_�1.�U��1��q�Q���8B�xv�,���%��e8�c�;&���hþ=�>���ǰ�E��4�)�=��X�SU�'8@����c5���Q�\��Hk����[/�4?��"�T�H�o0 ǡ������h+}n�L���^��N�:n}��#�:ːzJꟕ~&�U��~�P�:Q��Q`����>�ߺQ����!��UF�^L�P�3�t}�c�5Z�Z��>*�JxA�#�VOn[�:q��#/Ic���ؼ�3J�����T�i������Lw����o��"�K�����ۓ@��O�,_s�L�EZRR!�ʨ�ڿ5�����\.$3=]}�4����Ƨ�T\��Э^��6"�z����j���!o�Rynl�k�����x��J�!�䣦��h��<���~�ӆ���5���A\̅r=Nd��4j����"q��X�F��Zm�YR�!|�L%�<���p���{\��b�j���u���f�uX\iC�n���2��_�����n�w���
y���II�%�Y�>���@���#H{�sL�tMU'�r>NA0)�U����tH���aӒ����}�Ցȡ_>���gQ-����3�G�)���z<1'7p�<��?�sȔھ��m��h},
e��Xj�9����ġD`��3;�j�u�?9��^�t(�D��=g����-�_G�Tp����8��B\��g��������C�����_'䖫LW��w����y^�L��� ��Ɣ5%�3���� �xgo��$���%�6?��S0��a�`N��AgJ�ǧ�F��֤E�!�0m�}�}���/���+Ed灦:m��L�m�e";i��G�t�z����/����a!�px�o ב��|��Ѐ����q�*/ˇsp��̋'����%�o�/p�8�i���D��\�QI���-h;$6�d�}�/^8]2�7�D��<�D�7�(g����R*�0�}�\N��y�Os��NƆmq��� ��<�k��bN3�%�SUQ�� t��
y���Nǵ×m�1�H�y3u|�����������g�~^��)�m'_$O��k i�%��i<�('_=~gCBA^T���eJ�|��q�㮲�g��9&�����LHt��ym��oz*m�*�mYV%����\�� ��y��Z,��Ծ��bRV�3�y�,^L3:I���9m.£��[���kf��g���X��6d�9u�?�����K���;͑���C Q�٪�1muz�0e�M���k�\oKr�~(E{��객��3��3��F��	v3�?	ItQ� ��@]4�.��RA��2��_h�C#��Sw��%�4�`�(�NO��y�s/F��4	+���a7l#T�HI�t$Y��Cs��,����>�B&�ue1�`�\��T;W�#1t�0�)��'H*۩�����؈6|�����Jʠ�ac����s���\��H��b=o�(���n��q��ډZ(~j�+`[�HH�"uVY�zД1�=�$��oL�U�hS?S'�H�kH�0|��,\*�����J��2�d�)��:G���5e�n�l��L&ǒ_9N��Ubvy�c
�6p�O��\�p�T���]�D�4 t+� {�6t
�[�$���m� �WEܦ8��(����}n� 'r�?R�c��3,su��I)҆Rd QSՅ����� �� S��t��r�z�/0�s
UM������
�d��!�v�Cr�/�i�кZD��z�ޡHXl���d���A��u���~Y��5Ŀ0�SjV�9\y78I@J>ՇCV�j>R�\Wi��#����0Fa�@(>��0�O�ޯ�$���)�`���)'+N(�wvȐ�H���)J��͗6l^Ʉ��3�ә|aHr���6�1��<4��R'��U��!�*]O^���~e�h�������ġ�Gf�~0Et~M4��ًm��Z�� �,m�7Dzw�����$��7�����Lr�EW5!+(�J�b�YCk.�_�M��*�{�_�D��S��.�>8И�mta�#{�"�T0=.�w#]񕵚]��D�X܆I/Of���pnG"�:l�ژGN/~���O�3���>�+l/L�(0nGy+*_�����|��r�Fo���!w%�2�Kh���
B�y$jQUF�;eDf6�����~��C�8�m0�TpZ yID�;?s�	e��-^@�YM�m(�K7j��U@՘��R�7�?�|�n��^<(B�m�	W����:�$�
���mk�C� �_��beڄ�w����#�w�)L�7L�S
���2^�Pfxj�]�J
n2I��e�Y�w��5@Q��z[0�}޶������8v럒��xͨK�	��^<ǲe^�&�Wf�%��K�R���C*�@Y��r��B�Y+�H�Z���_��Y,u��L7B��i���<c��h�>m��������{ K��b�m���a��M2�(`�?�fK*W*J�y	d>�k��N�V�j��_���ʒKy���촷��ܜq��_����}�1R�jL���rJv=�
��(b'#���"���̇��Y`
������r��u�NKh��9k��%�$�ls(A�j�N�z��h@�T�)C�3~�dc��t��ҲY�����G�U,H,d��ξ?�83��j���V"w�^4�\N��6��,"+��v��]�qu��nS2����g��i�vt�<���'�Q�.�{n,������5BH���� �T}�`N{��s�%~Bwj%n��8�ܒ���=9�k���l��͍�T^j�(Z{�Q�	�X�$8����a����	 �P�E��}�{q$�[9����k�x,��8&7���՜��ӻ1���S�~��[��C����<���A?���,��p�Y��,�b֋�I	�.������dĽ�Fa�r�}�"�I�0c��'�mk�Ƃ`��������% �xЀ͖FͿ���e�Up�!�S�Y���2�M,�*5��%�⊧Ty������6� Ast���3��)J�~<)f���*^Z\&{�=��!�F$��KT�[%a!�y��}!�g^���?��zR`�zT�s�1�[Z򜬃GJ�n�+JΊ��oaִ����gk9'ρ$�O�jy�Ag2}j߸b��+�n�W�Ǉ�{�� �zdq�����[������:��+��~;���2Ck97(���S|��\M�ǦiW�'V�Σu�	V0ͥ�jɽ����$D�"q�j����(�޷�託�i��3�!Q�3�����fM)|@9NBPö��ͅX<��Y�� �7�҆G6��Ha�IP,W�&�b�Q[�C���M���8�$f�p�{L�\��\���申���*)�ȁ8X"J�3jRW��$��Ģ(�y�G�S�s��4�P��( ^p�2ش�A�z���#����x�+qg��A@��֛i�,���1��V(I�*-�!�r��.�?ս��sa��3��r�
�{kR��ph�sd�[��h'z���7�^&ɚJ�jÞ��6����̴Ì�